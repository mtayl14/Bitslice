* NGSPICE file created from bitslice.ext - technology: sky130A

.subckt inverter A B gnd vdd
X0 B A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X1 B A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
C0 A vdd 0.105f
C1 A B 0.0573f
C2 vdd B 0.0828f
C3 B gnd 0.32f
C4 A gnd 0.405f
C5 vdd gnd 0.456f
.ends

.subckt mux21 A B Y S gnd vdd S_n
X0 Y S A vdd sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X1 S_n S gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X2 B S Y gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 S_n S vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
X4 B S_n Y vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X5 Y S_n A gnd sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
C0 Y S_n 0.122f
C1 Y vdd 0.0197f
C2 Y A 0.175f
C3 Y S 0.12f
C4 Y B 0.175f
C5 S_n vdd 0.186f
C6 S_n A 0.232f
C7 S_n S 0.421f
C8 B S_n 0.101f
C9 A vdd 0.0531f
C10 S vdd 0.155f
C11 B vdd 0.0456f
C12 S A 0.101f
C13 B A 0.129f
C14 B S 0.0905f
C15 B gnd 0.249f
C16 Y gnd 0.11f
C17 A gnd 0.176f
C18 S gnd 0.621f
C19 vdd gnd 0.843f
C20 S_n gnd 0.433f
.ends

.subckt buffer_fo4 A B gnd vdd a_n240_0#
X0 a_n240_0# A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
X1 B a_n240_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.47 pd=3.92 as=0.504 ps=3.96 w=1.68 l=0.15
X2 a_n240_0# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X3 vdd a_n240_0# B vdd sky130_fd_pr__pfet_01v8 ad=1.01 pd=7.32 as=0.941 ps=7.28 w=3.36 l=0.15
C0 A vdd 0.118f
C1 A B 0.00714f
C2 a_n240_0# A 0.0759f
C3 B vdd 0.294f
C4 a_n240_0# vdd 0.267f
C5 a_n240_0# B 0.11f
C6 B gnd 0.415f
C7 A gnd 0.384f
C8 vdd gnd 1.67f
C9 a_n240_0# gnd 0.477f
.ends

.subckt addf A B CI gnd S CO vdd a_526_521# a_368_115# a_952_115# a_368_521# a_952_521#
+ a_784_115# a_27_115# a_27_521# CON a_870_115# a_870_521# a_526_115#
X0 a_952_521# CI a_870_521# vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.52 as=0.164 ps=1.52 w=1.26 l=0.15
X1 S a_784_115# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.334 pd=3.05 as=0.214 ps=1.6 w=1.26 l=0.15
X2 a_526_115# CI gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X3 a_27_521# B vdd vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X4 a_952_115# CI a_870_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0676 pd=0.78 as=0.0676 ps=0.78 w=0.52 l=0.15
X5 S a_784_115# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.57 as=0.0884 ps=0.86 w=0.52 l=0.15
X6 vdd A a_27_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.334 ps=3.05 w=1.26 l=0.15
X7 a_784_115# CON a_526_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X8 a_27_115# B gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X9 gnd A a_27_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.138 ps=1.57 w=0.52 l=0.15
X10 a_784_115# CON a_526_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X11 CON CI a_27_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X12 vdd A a_368_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.132 ps=1.47 w=1.26 l=0.15
X13 a_526_521# A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X14 CO CON vdd vdd sky130_fd_pr__pfet_01v8 ad=0.334 pd=3.05 as=0.334 ps=3.05 w=1.26 l=0.15
X15 CON CI a_27_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X16 a_870_521# B a_784_115# vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.52 as=0.176 ps=1.54 w=1.26 l=0.15
X17 gnd A a_368_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0546 ps=0.73 w=0.52 l=0.15
X18 a_526_115# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X19 CO CON gnd gnd sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.57 as=0.138 ps=1.57 w=0.52 l=0.15
X20 a_870_115# B a_784_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0676 pd=0.78 as=0.0728 ps=0.8 w=0.52 l=0.15
X21 a_368_521# B CON vdd sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.47 as=0.176 ps=1.54 w=1.26 l=0.15
X22 vdd B a_526_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X23 vdd A a_952_521# vdd sky130_fd_pr__pfet_01v8 ad=0.214 pd=1.6 as=0.164 ps=1.52 w=1.26 l=0.15
X24 a_368_115# B CON gnd sky130_fd_pr__nfet_01v8 ad=0.0546 pd=0.73 as=0.0728 ps=0.8 w=0.52 l=0.15
X25 gnd B a_526_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X26 gnd A a_952_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0884 pd=0.86 as=0.0676 ps=0.78 w=0.52 l=0.15
X27 a_526_521# CI vdd vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
C0 B a_870_521# 0.0013f
C1 B S 8.48e-19
C2 CON a_870_115# 0.00206f
C3 A S 0.0302f
C4 a_870_521# a_784_115# 0.0133f
C5 S a_784_115# 0.116f
C6 S CO 0.0234f
C7 CI a_870_521# 0.00263f
C8 B a_870_115# 2.05e-19
C9 CI S 0.00855f
C10 a_27_521# S 2.01e-19
C11 a_870_115# a_784_115# 0.00424f
C12 CON a_368_115# 0.00392f
C13 a_368_521# S 1.28e-19
C14 CON a_952_115# 0.0023f
C15 vdd a_368_115# 1.02e-19
C16 CON a_526_521# 0.00595f
C17 B a_368_115# 9.37e-19
C18 vdd a_526_521# 0.175f
C19 a_368_115# a_526_115# 6.28e-19
C20 B a_526_521# 0.036f
C21 A a_952_115# 3.88e-19
C22 vdd a_952_521# 0.00973f
C23 A a_526_521# 0.00216f
C24 a_952_115# a_784_115# 0.00282f
C25 CON vdd 0.165f
C26 a_526_521# a_526_115# 0.00723f
C27 a_526_521# a_784_115# 0.0546f
C28 A a_952_521# 0.00141f
C29 CI a_952_115# 5.65e-19
C30 B CON 0.28f
C31 CI a_526_521# 0.023f
C32 a_952_521# a_784_115# 0.0127f
C33 CON A 0.447f
C34 B vdd 0.294f
C35 CON a_526_115# 0.0472f
C36 a_870_521# S 7.59e-19
C37 CON a_784_115# 0.173f
C38 CI a_952_521# 0.00174f
C39 A vdd 0.169f
C40 CON CO 0.127f
C41 CON CI 0.219f
C42 vdd a_526_115# 0.00164f
C43 B A 0.511f
C44 vdd a_784_115# 0.149f
C45 CON a_27_521# 0.066f
C46 B a_526_115# 0.0263f
C47 vdd CO 0.11f
C48 B a_784_115# 0.19f
C49 vdd CI 0.122f
C50 a_870_115# S 3.84e-19
C51 A a_526_115# 0.00873f
C52 vdd a_27_521# 0.134f
C53 B CO 0.00429f
C54 A a_784_115# 0.19f
C55 a_368_521# CON 0.00367f
C56 B CI 0.88f
C57 B a_27_521# 0.0591f
C58 a_784_115# a_526_115# 0.0359f
C59 A CO 7.16e-19
C60 A CI 0.503f
C61 a_368_521# vdd 0.00893f
C62 A a_27_521# 0.0145f
C63 CO a_784_115# 0.00108f
C64 CI a_526_115# 0.0258f
C65 CI a_784_115# 0.0932f
C66 CON a_27_115# 0.05f
C67 a_368_521# B 0.00709f
C68 CI CO 4.26e-19
C69 vdd a_27_115# 8.57e-19
C70 CI a_27_521# 0.00307f
C71 a_368_521# a_784_115# 5.73e-19
C72 B a_27_115# 0.0277f
C73 a_952_115# S 7.1e-19
C74 A a_27_115# 0.0471f
C75 a_526_521# S 6.86e-19
C76 a_952_521# S 0.00114f
C77 CI a_27_115# 0.00565f
C78 a_27_115# a_27_521# 0.00483f
C79 CON S 0.113f
C80 vdd a_870_521# 0.00633f
C81 vdd S 0.139f
C82 CO gnd 0.209f
C83 S gnd 0.116f
C84 CI gnd 0.525f
C85 B gnd 0.705f
C86 A gnd 0.804f
C87 vdd gnd 2.33f
C88 a_952_115# gnd 0.00647f
C89 a_870_115# gnd 0.00354f
C90 a_526_115# gnd 0.155f
C91 a_368_115# gnd 0.00506f
C92 a_27_115# gnd 0.159f
C93 a_952_521# gnd 1.04e-19
C94 a_870_521# gnd 9.72e-21
C95 a_526_521# gnd 0.0201f
C96 a_368_521# gnd 2.66e-19
C97 a_27_521# gnd 0.057f
C98 a_784_115# gnd 0.291f
C99 CON gnd 0.802f
.ends

.subckt d_flip_flop CLK D Q gnd vdd a_494_0# a_1248_0# CLK_n a_220_426# a_494_426#
+ a_974_426# a_220_0# inverter_1_out common_2 common_1 a_974_0# a_1248_426#
X0 inverter_1_out common_1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X1 gnd inverter_1_out a_494_0# gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
X2 common_2 CLK_n a_974_426# vdd sky130_fd_pr__pfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 gnd Q a_1248_0# gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
X4 a_974_0# inverter_1_out gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X5 a_220_426# D vdd vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X6 a_494_0# CLK common_1 gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X7 a_1248_0# CLK_n common_2 gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X8 CLK_n CLK vdd vdd sky130_fd_pr__pfet_01v8 ad=0.445 pd=3.89 as=0.445 ps=3.89 w=1.68 l=0.15
X9 common_1 CLK a_220_426# vdd sky130_fd_pr__pfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X10 Q common_2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.34 pd=2.8 as=0.134 ps=1.23 w=0.84 l=0.15
X11 a_1248_426# CLK common_2 vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X12 CLK_n CLK gnd gnd sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
X13 common_1 CLK_n a_220_0# gnd sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X14 vdd Q a_1248_426# vdd sky130_fd_pr__pfet_01v8 ad=0.134 pd=1.23 as=0.0819 ps=0.81 w=0.42 l=0.15
X15 common_2 CLK a_974_0# gnd sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X16 inverter_1_out common_1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X17 Q common_2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X18 a_494_426# CLK_n common_1 vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X19 a_974_426# inverter_1_out vdd vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X20 a_220_0# D gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X21 vdd inverter_1_out a_494_426# vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
C0 common_1 D 0.0338f
C1 a_220_0# CLK 0.00497f
C2 a_494_0# vdd 2.34e-19
C3 common_1 CLK 0.294f
C4 D CLK_n 0.122f
C5 vdd a_220_426# 0.00638f
C6 CLK_n CLK 1.39f
C7 a_1248_0# CLK_n 0.00313f
C8 inverter_1_out common_2 0.0217f
C9 D CLK 0.188f
C10 a_494_0# Q 1.34e-19
C11 vdd common_2 0.165f
C12 common_1 inverter_1_out 0.241f
C13 common_1 vdd 0.175f
C14 CLK_n inverter_1_out 0.21f
C15 vdd CLK_n 0.318f
C16 D inverter_1_out 0.00602f
C17 Q common_2 0.269f
C18 inverter_1_out CLK 0.224f
C19 D vdd 0.109f
C20 a_1248_426# common_2 0.00273f
C21 a_220_0# Q 1.24e-19
C22 vdd CLK 0.661f
C23 a_1248_0# vdd 3.63e-19
C24 Q common_1 2.17e-19
C25 a_974_0# common_2 0.00277f
C26 Q CLK_n 0.0719f
C27 Q D 2.13e-19
C28 Q CLK 0.0622f
C29 Q a_1248_0# 9.54e-19
C30 vdd inverter_1_out 0.302f
C31 a_974_0# CLK_n 0.00401f
C32 a_974_426# common_2 0.00211f
C33 CLK a_1248_426# 0.0028f
C34 a_974_0# CLK 0.00228f
C35 common_1 a_494_426# 0.00211f
C36 a_494_0# common_2 2.69e-19
C37 a_974_426# CLK_n 0.00166f
C38 Q inverter_1_out 0.00505f
C39 Q vdd 0.172f
C40 a_494_426# CLK_n 0.00166f
C41 vdd a_1248_426# 0.00627f
C42 a_974_426# CLK 0.00292f
C43 a_494_426# CLK 0.00292f
C44 a_494_0# CLK_n 0.00356f
C45 a_974_0# vdd 2.34e-19
C46 common_1 a_220_426# 0.00211f
C47 a_220_0# common_2 9.78e-20
C48 a_494_0# CLK 0.00903f
C49 common_1 common_2 3.81e-19
C50 CLK_n a_220_426# 6.84e-19
C51 a_220_0# common_1 0.00135f
C52 a_974_426# vdd 0.00744f
C53 Q a_974_0# 3.81e-19
C54 CLK a_220_426# 0.00458f
C55 CLK_n common_2 0.209f
C56 D common_2 1.9e-19
C57 a_494_426# vdd 0.00747f
C58 a_220_0# CLK_n 0.00636f
C59 common_1 CLK_n 0.257f
C60 CLK common_2 0.116f
C61 a_1248_0# common_2 0.00945f
C62 Q gnd 0.492f
C63 D gnd 0.27f
C64 CLK gnd 1.15f
C65 vdd gnd 2.63f
C66 a_1248_0# gnd 0.00421f
C67 a_974_0# gnd 0.00647f
C68 a_494_0# gnd 0.00449f
C69 a_220_0# gnd 0.00356f
C70 a_1248_426# gnd 2.68e-19
C71 a_974_426# gnd 2.68e-19
C72 a_494_426# gnd 2.68e-19
C73 common_2 gnd 0.517f
C74 common_1 gnd 0.302f
C75 inverter_1_out gnd 0.593f
C76 CLK_n gnd 0.855f
.ends

.subckt and2 A B Y gnd vdd a_30_n42# Y_n
X0 vdd B Y_n vdd sky130_fd_pr__pfet_01v8 ad=0.212 pd=1.35 as=0.118 ps=1.12 w=0.84 l=0.15
X1 Y Y_n vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.212 ps=1.35 w=0.84 l=0.15
X2 Y Y_n gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.159 ps=1.35 w=0.42 l=0.15
X3 Y_n A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X4 gnd B a_30_n42# gnd sky130_fd_pr__nfet_01v8 ad=0.159 pd=1.35 as=0.118 ps=1.12 w=0.84 l=0.15
X5 a_30_n42# A Y_n gnd sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
C0 vdd a_30_n42# 4.51e-19
C1 a_30_n42# Y 9.31e-19
C2 B A 0.0938f
C3 Y_n a_30_n42# 0.0116f
C4 vdd A 0.072f
C5 vdd B 0.108f
C6 A Y 0.00134f
C7 B Y 0.0233f
C8 vdd Y 0.0836f
C9 A Y_n 0.0914f
C10 B Y_n 0.176f
C11 vdd Y_n 0.186f
C12 Y_n Y 0.0794f
C13 Y gnd 0.284f
C14 B gnd 0.248f
C15 A gnd 0.322f
C16 vdd gnd 0.757f
C17 a_30_n42# gnd 0.00713f
C18 Y_n gnd 0.444f
.ends

.subckt register D CLK EN Q vdd d_flip_flop_0/a_494_426# d_flip_flop_0/a_974_426#
+ and2_0/Y_n d_flip_flop_0/common_2 d_flip_flop_0/common_1 and2_0/Y d_flip_flop_0/a_974_0#
+ d_flip_flop_0/a_1248_426# d_flip_flop_0/a_494_0# and2_0/a_30_n42# d_flip_flop_0/inverter_1_out
+ d_flip_flop_0/a_1248_0# d_flip_flop_0/CLK_n gnd d_flip_flop_0/a_220_426#
Xd_flip_flop_0 and2_0/Y D Q gnd vdd d_flip_flop_0/a_494_0# d_flip_flop_0/a_1248_0#
+ d_flip_flop_0/CLK_n d_flip_flop_0/a_220_426# d_flip_flop_0/a_494_426# d_flip_flop_0/a_974_426#
+ d_flip_flop_0/a_220_0# d_flip_flop_0/inverter_1_out d_flip_flop_0/common_2 d_flip_flop_0/common_1
+ d_flip_flop_0/a_974_0# d_flip_flop_0/a_1248_426# d_flip_flop
Xand2_0 CLK EN and2_0/Y gnd vdd and2_0/a_30_n42# and2_0/Y_n and2
C0 CLK D 4.88e-20
C1 EN d_flip_flop_0/common_1 2.23e-19
C2 CLK and2_0/Y 0.0199f
C3 and2_0/Y D 0.00132f
C4 vdd D 0.00388f
C5 CLK and2_0/Y_n 2.84e-32
C6 d_flip_flop_0/a_1248_0# and2_0/Y 8.55e-20
C7 Q and2_0/Y 1.66e-19
C8 and2_0/Y_n D 0.00817f
C9 vdd and2_0/Y 0.0522f
C10 and2_0/Y_n and2_0/Y 0.0383f
C11 vdd and2_0/Y_n 0.014f
C12 EN CLK -1.42e-32
C13 EN D 7.78e-19
C14 EN Q 2.99e-20
C15 EN and2_0/Y 0.0186f
C16 vdd EN 0.00216f
C17 and2_0/Y d_flip_flop_0/CLK_n 0.0351f
C18 vdd d_flip_flop_0/CLK_n 5.37e-19
C19 d_flip_flop_0/inverter_1_out and2_0/Y 7.03e-19
C20 and2_0/Y_n d_flip_flop_0/CLK_n 5.91e-19
C21 and2_0/Y d_flip_flop_0/common_2 3.33e-19
C22 Q d_flip_flop_0/a_220_0# -1.39e-35
C23 and2_0/Y d_flip_flop_0/a_974_0# 1.25e-19
C24 and2_0/Y d_flip_flop_0/a_220_0# 6.81e-19
C25 EN d_flip_flop_0/CLK_n 0.00102f
C26 d_flip_flop_0/inverter_1_out EN 1.44e-19
C27 EN d_flip_flop_0/common_2 3.89e-20
C28 and2_0/Y d_flip_flop_0/common_1 9.82e-19
C29 and2_0/Y d_flip_flop_0/a_494_0# 2.46e-19
C30 and2_0/a_30_n42# and2_0/Y 7.24e-19
C31 vdd gnd 3.28f
C32 EN gnd 0.231f
C33 CLK gnd 0.306f
C34 and2_0/a_30_n42# gnd 0.00713f
C35 and2_0/Y_n gnd 0.445f
C36 Q gnd 0.492f
C37 D gnd 0.257f
C38 and2_0/Y gnd 1.29f
C39 d_flip_flop_0/a_1248_0# gnd 0.00421f
C40 d_flip_flop_0/a_974_0# gnd 0.00647f
C41 d_flip_flop_0/a_494_0# gnd 0.00449f
C42 d_flip_flop_0/a_220_0# gnd 0.00356f
C43 d_flip_flop_0/a_1248_426# gnd 2.68e-19
C44 d_flip_flop_0/a_974_426# gnd 2.68e-19
C45 d_flip_flop_0/a_494_426# gnd 2.68e-19
C46 d_flip_flop_0/common_2 gnd 0.517f
C47 d_flip_flop_0/common_1 gnd 0.302f
C48 d_flip_flop_0/inverter_1_out gnd 0.593f
C49 d_flip_flop_0/CLK_n gnd 0.855f
.ends

.subckt bitslice gnd vdd B A SUB CI STORE CLK CO Q
Xinverter_0 B mux21_0/B gnd vdd inverter
Xmux21_0 B mux21_0/B addf_0/B SUB gnd vdd mux21_0/S_n mux21
Xbuffer_fo4_0 CLK register_0/CLK gnd vdd buffer_fo4_0/a_n240_0# buffer_fo4
Xaddf_0 A addf_0/B CI gnd addf_0/S CO vdd addf_0/a_526_521# addf_0/a_368_115# addf_0/a_952_115#
+ addf_0/a_368_521# addf_0/a_952_521# addf_0/a_784_115# addf_0/a_27_115# addf_0/a_27_521#
+ addf_0/CON addf_0/a_870_115# addf_0/a_870_521# addf_0/a_526_115# addf
Xregister_0 addf_0/S register_0/CLK STORE Q vdd register_0/d_flip_flop_0/a_494_426#
+ register_0/d_flip_flop_0/a_974_426# register_0/and2_0/Y_n register_0/d_flip_flop_0/common_2
+ register_0/d_flip_flop_0/common_1 register_0/and2_0/Y register_0/d_flip_flop_0/a_974_0#
+ register_0/d_flip_flop_0/a_1248_426# register_0/d_flip_flop_0/a_494_0# register_0/and2_0/a_30_n42#
+ register_0/d_flip_flop_0/inverter_1_out register_0/d_flip_flop_0/a_1248_0# register_0/d_flip_flop_0/CLK_n
+ gnd register_0/d_flip_flop_0/a_220_426# register
C0 A addf_0/B 0.138f
C1 addf_0/a_368_521# addf_0/B 0.00251f
C2 addf_0/a_952_115# mux21_0/B 1.85e-19
C3 addf_0/a_870_115# mux21_0/B 1.93e-19
C4 addf_0/S vdd 0.988f
C5 register_0/d_flip_flop_0/common_1 buffer_fo4_0/a_n240_0# 1.91e-20
C6 mux21_0/B addf_0/a_526_115# 6.04e-19
C7 addf_0/a_27_521# addf_0/CON 1.42e-32
C8 mux21_0/B addf_0/a_784_115# 3.13e-19
C9 SUB vdd 0.0757f
C10 STORE vdd 0.101f
C11 addf_0/a_27_521# CO 0.0063f
C12 buffer_fo4_0/a_n240_0# addf_0/CON 0.00294f
C13 addf_0/B addf_0/a_784_115# 0.00117f
C14 register_0/CLK vdd -0.0106f
C15 register_0/d_flip_flop_0/inverter_1_out buffer_fo4_0/a_n240_0# 9.01e-21
C16 CI addf_0/a_27_115# 0.0106f
C17 mux21_0/S_n addf_0/CON 6.69e-19
C18 CI addf_0/a_27_521# 0.00157f
C19 addf_0/a_870_521# addf_0/B 6.35e-19
C20 CLK vdd 0.113f
C21 register_0/d_flip_flop_0/CLK_n buffer_fo4_0/a_n240_0# 1.5e-19
C22 buffer_fo4_0/a_n240_0# CO 0.0328f
C23 addf_0/B mux21_0/B 0.114f
C24 B vdd -0.026f
C25 addf_0/a_952_521# addf_0/B 5.33e-19
C26 mux21_0/S_n CO 6.34e-19
C27 register_0/and2_0/a_30_n42# vdd -4.51e-19
C28 addf_0/S SUB 9.42e-21
C29 CI buffer_fo4_0/a_n240_0# 2.83e-19
C30 register_0/and2_0/Y_n vdd -0.00765f
C31 A addf_0/a_27_115# 0.00248f
C32 addf_0/S STORE 0.115f
C33 CI mux21_0/S_n 4.53e-19
C34 register_0/and2_0/Y vdd -0.0125f
C35 A addf_0/a_27_521# 0.0163f
C36 buffer_fo4_0/a_n240_0# addf_0/a_526_521# 4.17e-21
C37 addf_0/S register_0/CLK 0.114f
C38 mux21_0/S_n addf_0/a_526_521# 3.39e-20
C39 addf_0/S CLK 0.0844f
C40 A buffer_fo4_0/a_n240_0# 4.29e-19
C41 addf_0/S register_0/and2_0/a_30_n42# 6.46e-19
C42 A mux21_0/S_n 0.0628f
C43 addf_0/S register_0/and2_0/Y_n 0.0285f
C44 addf_0/S Q 8.38e-19
C45 STORE register_0/CLK 0.0421f
C46 addf_0/S register_0/and2_0/Y 0.133f
C47 CLK SUB 3.14e-19
C48 STORE CLK 0.0414f
C49 SUB B 0.312f
C50 CLK register_0/CLK 0.0245f
C51 STORE register_0/and2_0/a_30_n42# 0.00131f
C52 STORE register_0/and2_0/Y_n 0.0262f
C53 STORE Q -4.62e-21
C54 register_0/CLK register_0/and2_0/a_30_n42# 9.08e-20
C55 buffer_fo4_0/a_n240_0# addf_0/a_526_115# 1.23e-20
C56 register_0/CLK register_0/and2_0/Y_n 0.0204f
C57 STORE register_0/and2_0/Y 0.0981f
C58 CLK register_0/and2_0/a_30_n42# 2.23e-19
C59 addf_0/S register_0/d_flip_flop_0/a_1248_426# 3.05e-19
C60 register_0/CLK register_0/and2_0/Y -0.00576f
C61 mux21_0/B addf_0/a_27_115# 0.039f
C62 CLK register_0/and2_0/Y_n 0.00172f
C63 addf_0/S register_0/d_flip_flop_0/a_974_426# 4.8e-19
C64 mux21_0/B addf_0/a_27_521# 0.0438f
C65 buffer_fo4_0/a_n240_0# addf_0/a_784_115# 1.9e-19
C66 STORE register_0/d_flip_flop_0/a_1248_0# 1.81e-20
C67 CLK register_0/and2_0/Y 2.23e-19
C68 addf_0/S register_0/d_flip_flop_0/a_494_426# 0.00125f
C69 register_0/d_flip_flop_0/a_974_0# STORE 2.57e-20
C70 mux21_0/S_n addf_0/a_784_115# 6.68e-20
C71 addf_0/B addf_0/a_27_115# 3.14e-19
C72 addf_0/S register_0/d_flip_flop_0/a_220_426# 0.00193f
C73 addf_0/CON vdd -0.00395f
C74 addf_0/B addf_0/a_27_521# 0.0554f
C75 register_0/and2_0/Y register_0/and2_0/a_30_n42# -4.89e-19
C76 register_0/d_flip_flop_0/a_494_0# STORE 3.46e-20
C77 addf_0/S register_0/d_flip_flop_0/common_2 0.0011f
C78 mux21_0/B buffer_fo4_0/a_n240_0# 2.44e-20
C79 register_0/and2_0/Y_n register_0/and2_0/Y -0.00662f
C80 addf_0/S register_0/d_flip_flop_0/common_1 0.00644f
C81 mux21_0/S_n mux21_0/B 0.0772f
C82 CO vdd 0.221f
C83 addf_0/B buffer_fo4_0/a_n240_0# 4.31e-20
C84 mux21_0/S_n addf_0/B 0.0787f
C85 CI vdd 2.71e-19
C86 STORE register_0/d_flip_flop_0/common_2 -1.32e-20
C87 addf_0/S addf_0/CON 0.0179f
C88 STORE register_0/d_flip_flop_0/common_1 -1.22e-19
C89 addf_0/S register_0/d_flip_flop_0/inverter_1_out 0.00305f
C90 register_0/d_flip_flop_0/CLK_n addf_0/S 0.0208f
C91 addf_0/S CO 0.0948f
C92 A vdd 0.347f
C93 CLK addf_0/a_368_115# 2.05e-19
C94 SUB addf_0/CON 0.00238f
C95 addf_0/S CI 0.00206f
C96 STORE addf_0/CON 4.04e-20
C97 STORE register_0/d_flip_flop_0/inverter_1_out 9.42e-20
C98 addf_0/S addf_0/a_526_521# 0.0015f
C99 register_0/CLK addf_0/CON 9.99e-19
C100 SUB CO 0.0126f
C101 register_0/d_flip_flop_0/CLK_n STORE 0.00234f
C102 STORE CO 1.05e-20
C103 CLK addf_0/CON 0.0414f
C104 register_0/CLK CO 2.92e-19
C105 CI SUB 0.0263f
C106 A addf_0/S 0.0025f
C107 B addf_0/CON 0.00295f
C108 register_0/and2_0/a_30_n42# addf_0/CON 2.07e-20
C109 register_0/and2_0/Y_n addf_0/CON 9.36e-20
C110 CLK CO 0.208f
C111 CI register_0/CLK 0.00174f
C112 addf_0/S addf_0/a_368_521# 3.02e-19
C113 register_0/and2_0/Y addf_0/CON 1.35e-19
C114 buffer_fo4_0/a_n240_0# addf_0/a_27_115# 1.58e-21
C115 CI CLK 0.0161f
C116 register_0/and2_0/Y_n CO 7.68e-21
C117 A SUB 0.181f
C118 addf_0/a_784_115# vdd -2.84e-32
C119 buffer_fo4_0/a_n240_0# addf_0/a_27_521# 3.21e-20
C120 CI B 3.54e-19
C121 CLK addf_0/a_526_521# 5.44e-19
C122 A STORE 2.4e-21
C123 register_0/and2_0/Y CO 3.66e-19
C124 mux21_0/S_n addf_0/a_27_521# 0.00253f
C125 A register_0/CLK 0.00152f
C126 mux21_0/B vdd 7.82e-19
C127 A CLK 0.00334f
C128 A B 0.139f
C129 addf_0/B vdd 0.174f
C130 addf_0/a_368_521# CLK 1.4e-19
C131 addf_0/S addf_0/a_784_115# 0.00572f
C132 A register_0/and2_0/Y_n 9.67e-21
C133 SUB addf_0/a_526_115# 3.39e-20
C134 addf_0/a_870_521# addf_0/S 0.00164f
C135 addf_0/S mux21_0/B 8.81e-20
C136 CLK addf_0/a_952_115# 7.72e-19
C137 addf_0/S addf_0/a_952_521# 0.00216f
C138 addf_0/a_870_115# CLK 5.86e-19
C139 SUB addf_0/a_784_115# 3.28e-20
C140 CLK addf_0/a_526_115# 0.00107f
C141 addf_0/S addf_0/B 0.00812f
C142 addf_0/a_368_115# CO 5.7e-19
C143 register_0/CLK addf_0/a_784_115# 9.51e-20
C144 SUB mux21_0/B 0.122f
C145 CLK addf_0/a_784_115# 0.00431f
C146 CI addf_0/a_368_115# 0.00109f
C147 SUB addf_0/B 0.00425f
C148 addf_0/a_870_521# CLK 4.45e-19
C149 CO addf_0/CON 0.105f
C150 CLK mux21_0/B 7.27e-20
C151 addf_0/a_952_521# CLK 6.32e-19
C152 register_0/CLK addf_0/B 2.48e-20
C153 addf_0/a_784_115# register_0/and2_0/Y 3.88e-21
C154 B mux21_0/B 0.154f
C155 CI addf_0/CON 0.027f
C156 CLK addf_0/B 0.00152f
C157 B addf_0/B 0.00835f
C158 addf_0/a_27_115# vdd -2.4e-19
C159 CI CO 0.0793f
C160 addf_0/a_27_521# vdd -0.00326f
C161 addf_0/a_526_521# CO 0.0216f
C162 A addf_0/CON 0.00319f
C163 buffer_fo4_0/a_n240_0# vdd -0.00691f
C164 mux21_0/S_n vdd -0.0175f
C165 A CO 0.125f
C166 addf_0/S addf_0/a_27_521# 1.38e-19
C167 A CI 0.0985f
C168 addf_0/a_368_521# CO 0.00464f
C169 A addf_0/a_526_521# 0.002f
C170 addf_0/S buffer_fo4_0/a_n240_0# 0.0578f
C171 SUB addf_0/a_27_115# 0.001f
C172 addf_0/a_952_115# CO 0.00134f
C173 addf_0/a_870_115# CO 6.29e-19
C174 addf_0/S mux21_0/S_n 1.96e-20
C175 SUB addf_0/a_27_521# 1.14e-21
C176 addf_0/a_368_115# mux21_0/B 6.27e-19
C177 addf_0/a_526_115# CO 0.00227f
C178 CI addf_0/a_952_115# 4.54e-19
C179 addf_0/a_870_115# CI 4.76e-19
C180 A addf_0/a_368_521# 0.00106f
C181 CLK addf_0/a_27_115# 9.61e-21
C182 SUB buffer_fo4_0/a_n240_0# 6.83e-22
C183 CI addf_0/a_526_115# 0.0032f
C184 CLK addf_0/a_27_521# 9.61e-21
C185 STORE buffer_fo4_0/a_n240_0# 0.00654f
C186 mux21_0/S_n SUB 0.0189f
C187 addf_0/a_784_115# CO 0.0517f
C188 B addf_0/a_27_115# 9.82e-20
C189 mux21_0/B addf_0/CON 0.00811f
C190 register_0/CLK buffer_fo4_0/a_n240_0# 0.00381f
C191 addf_0/a_870_521# CO 0.00527f
C192 CI addf_0/a_784_115# 0.00184f
C193 addf_0/B addf_0/CON 0.00968f
C194 CLK buffer_fo4_0/a_n240_0# 0.0335f
C195 mux21_0/B CO 6.7e-20
C196 addf_0/a_952_521# CO 0.00514f
C197 mux21_0/S_n CLK 6.71e-19
C198 mux21_0/S_n B 0.0591f
C199 CI mux21_0/B 0.0259f
C200 addf_0/B CO 0.0652f
C201 buffer_fo4_0/a_n240_0# register_0/and2_0/Y_n 0.00291f
C202 buffer_fo4_0/a_n240_0# register_0/and2_0/Y 0.00145f
C203 A addf_0/a_784_115# 0.00104f
C204 CI addf_0/B 0.031f
C205 A addf_0/a_870_521# 3.54e-19
C206 addf_0/B addf_0/a_526_521# 0.00279f
C207 A mux21_0/B 0.194f
C208 vdd gnd 8.03f
C209 addf_0/S gnd 0.564f
C210 STORE gnd 0.398f
C211 register_0/CLK gnd 0.66f
C212 register_0/and2_0/a_30_n42# gnd 0.00755f
C213 register_0/and2_0/Y_n gnd 0.448f
C214 Q gnd 0.492f
C215 register_0/and2_0/Y gnd 1.26f
C216 register_0/d_flip_flop_0/a_1248_0# gnd 0.00421f
C217 register_0/d_flip_flop_0/a_974_0# gnd 0.00647f
C218 register_0/d_flip_flop_0/a_494_0# gnd 0.00449f
C219 register_0/d_flip_flop_0/a_220_0# gnd 0.00356f
C220 register_0/d_flip_flop_0/a_1248_426# gnd 2.68e-19
C221 register_0/d_flip_flop_0/a_974_426# gnd 2.68e-19
C222 register_0/d_flip_flop_0/a_494_426# gnd 2.68e-19
C223 register_0/d_flip_flop_0/common_2 gnd 0.517f
C224 register_0/d_flip_flop_0/common_1 gnd 0.302f
C225 register_0/d_flip_flop_0/inverter_1_out gnd 0.593f
C226 register_0/d_flip_flop_0/CLK_n gnd 0.855f
C227 CO gnd 0.466f
C228 CI gnd 0.635f
C229 A gnd 0.941f
C230 addf_0/a_952_115# gnd 0.00647f
C231 addf_0/a_870_115# gnd 0.00354f
C232 addf_0/a_526_115# gnd 0.155f
C233 addf_0/a_368_115# gnd 0.00506f
C234 addf_0/a_27_115# gnd 0.162f
C235 addf_0/a_952_521# gnd 1.04e-19
C236 addf_0/a_870_521# gnd 9.72e-21
C237 addf_0/a_526_521# gnd 0.0201f
C238 addf_0/a_368_521# gnd 2.66e-19
C239 addf_0/a_27_521# gnd 0.0569f
C240 addf_0/a_784_115# gnd 0.291f
C241 addf_0/CON gnd 0.804f
C242 CLK gnd 0.463f
C243 buffer_fo4_0/a_n240_0# gnd 0.476f
C244 mux21_0/B gnd 0.644f
C245 addf_0/B gnd 0.766f
C246 B gnd 0.484f
C247 SUB gnd 0.718f
C248 mux21_0/S_n gnd 0.413f
.ends

