* NGSPICE file created from and2.ext - technology: sky130A

.subckt and2 A B Y
X0 w_n98_348# B Y_n w_n98_348# sky130_fd_pr__pfet_01v8 ad=0.212 pd=1.35 as=0.118 ps=1.12 w=0.84 l=0.15
X1 Y Y_n w_n98_348# w_n98_348# sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.212 ps=1.35 w=0.84 l=0.15
X2 Y Y_n a_n2_n145# a_n2_n145# sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.159 ps=1.35 w=0.42 l=0.15
X3 Y_n A w_n98_348# w_n98_348# sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X4 a_n2_n145# B a_30_n42# a_n2_n145# sky130_fd_pr__nfet_01v8 ad=0.159 pd=1.35 as=0.118 ps=1.12 w=0.84 l=0.15
X5 a_30_n42# A Y_n a_n2_n145# sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
.ends

