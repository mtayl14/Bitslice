magic
tech sky130A
magscale 1 2
timestamp 1701814136
<< nwell >>
rect -98 348 1612 706
rect -98 264 119 348
<< nmos >>
rect 0 -42 30 126
rect 190 0 220 84
rect 298 0 328 84
rect 464 0 494 84
rect 572 0 602 84
rect 680 0 710 84
rect 944 0 974 84
rect 1052 0 1082 84
rect 1218 0 1248 84
rect 1326 0 1356 84
rect 1434 0 1464 84
<< pmos >>
rect 0 300 30 636
rect 190 426 220 510
rect 298 426 328 510
rect 464 426 494 510
rect 572 426 602 510
rect 680 426 710 510
rect 944 426 974 510
rect 1052 426 1082 510
rect 1218 426 1248 510
rect 1326 426 1356 510
rect 1434 384 1464 552
<< ndiff >>
rect -53 68 0 126
rect -53 16 -45 68
rect -11 16 0 68
rect -53 -42 0 16
rect 30 68 83 126
rect 30 16 41 68
rect 75 16 83 68
rect 30 -42 83 16
rect 137 68 190 84
rect 137 16 145 68
rect 179 16 190 68
rect 137 0 190 16
rect 220 0 298 84
rect 328 68 464 84
rect 328 16 379 68
rect 413 16 464 68
rect 328 0 464 16
rect 494 0 572 84
rect 602 68 680 84
rect 602 16 624 68
rect 658 16 680 68
rect 602 0 680 16
rect 710 68 822 84
rect 710 16 780 68
rect 814 16 822 68
rect 710 0 822 16
rect 891 68 944 84
rect 891 16 899 68
rect 933 16 944 68
rect 891 0 944 16
rect 974 0 1052 84
rect 1082 68 1218 84
rect 1082 16 1133 68
rect 1167 16 1218 68
rect 1082 0 1218 16
rect 1248 0 1326 84
rect 1356 68 1434 84
rect 1356 16 1378 68
rect 1412 16 1434 68
rect 1356 0 1434 16
rect 1464 68 1576 84
rect 1464 16 1534 68
rect 1568 16 1576 68
rect 1464 0 1576 16
<< pdiff >>
rect -53 536 0 636
rect -53 400 -45 536
rect -11 400 0 536
rect -53 300 0 400
rect 30 536 83 636
rect 30 400 41 536
rect 75 400 83 536
rect 1384 510 1434 552
rect 137 492 190 510
rect 137 458 145 492
rect 179 458 190 492
rect 137 426 190 458
rect 220 426 298 510
rect 328 494 464 510
rect 328 460 379 494
rect 413 460 464 494
rect 328 426 464 460
rect 494 426 572 510
rect 602 494 680 510
rect 602 460 624 494
rect 658 460 680 494
rect 602 426 680 460
rect 710 494 822 510
rect 710 460 780 494
rect 814 460 822 494
rect 710 426 822 460
rect 891 494 944 510
rect 891 460 899 494
rect 933 460 944 494
rect 891 426 944 460
rect 974 426 1052 510
rect 1082 494 1218 510
rect 1082 460 1133 494
rect 1167 460 1218 494
rect 1082 426 1218 460
rect 1248 426 1326 510
rect 1356 494 1434 510
rect 1356 460 1378 494
rect 1412 460 1434 494
rect 1356 426 1434 460
rect 30 300 83 400
rect 1384 384 1434 426
rect 1464 510 1514 552
rect 1464 494 1576 510
rect 1464 460 1534 494
rect 1568 460 1576 494
rect 1464 426 1576 460
rect 1464 384 1514 426
<< ndiffc >>
rect -45 16 -11 68
rect 41 16 75 68
rect 145 16 179 68
rect 379 16 413 68
rect 624 16 658 68
rect 780 16 814 68
rect 899 16 933 68
rect 1133 16 1167 68
rect 1378 16 1412 68
rect 1534 16 1568 68
<< pdiffc >>
rect -45 400 -11 536
rect 41 400 75 536
rect 145 458 179 492
rect 379 460 413 494
rect 624 460 658 494
rect 780 460 814 494
rect 899 460 933 494
rect 1133 460 1167 494
rect 1378 460 1412 494
rect 1534 460 1568 494
<< psubdiff >>
rect 23 -145 48 -111
rect 82 -145 107 -111
rect 223 -118 248 -84
rect 282 -118 307 -84
rect 423 -118 448 -84
rect 482 -118 507 -84
rect 623 -118 648 -84
rect 682 -118 707 -84
rect 823 -118 848 -84
rect 882 -118 907 -84
rect 1023 -118 1048 -84
rect 1082 -118 1107 -84
rect 1223 -118 1248 -84
rect 1282 -118 1307 -84
rect 1423 -118 1448 -84
rect 1482 -118 1507 -84
<< nsubdiff >>
rect 223 636 248 670
rect 282 636 307 670
rect 423 636 448 670
rect 482 636 507 670
rect 623 636 648 670
rect 682 636 707 670
rect 823 636 848 670
rect 882 636 907 670
rect 1023 636 1048 670
rect 1082 636 1107 670
rect 1223 636 1248 670
rect 1282 636 1307 670
rect 1423 636 1448 670
rect 1482 636 1507 670
<< psubdiffcont >>
rect 48 -145 82 -111
rect 248 -118 282 -84
rect 448 -118 482 -84
rect 648 -118 682 -84
rect 848 -118 882 -84
rect 1048 -118 1082 -84
rect 1248 -118 1282 -84
rect 1448 -118 1482 -84
<< nsubdiffcont >>
rect 248 636 282 670
rect 448 636 482 670
rect 648 636 682 670
rect 848 636 882 670
rect 1048 636 1082 670
rect 1248 636 1282 670
rect 1448 636 1482 670
<< poly >>
rect 0 636 30 666
rect 190 510 220 582
rect 298 510 328 582
rect 464 510 494 582
rect 572 510 602 582
rect 680 510 710 582
rect 944 510 974 582
rect 1052 510 1082 582
rect 1218 510 1248 582
rect 1326 510 1356 582
rect 1434 552 1464 582
rect 0 266 30 300
rect -66 250 30 266
rect 190 252 220 426
rect 298 350 328 426
rect 262 334 328 350
rect 262 300 278 334
rect 312 300 328 334
rect 262 284 328 300
rect 464 350 494 426
rect 464 334 530 350
rect 464 300 480 334
rect 514 300 530 334
rect 464 284 530 300
rect -66 216 -50 250
rect -16 216 30 250
rect -66 200 30 216
rect 0 126 30 200
rect 154 236 220 252
rect 154 202 170 236
rect 204 202 220 236
rect 154 186 220 202
rect 190 84 220 186
rect 572 184 602 426
rect 680 290 710 426
rect 662 274 728 290
rect 662 240 678 274
rect 712 240 728 274
rect 944 250 974 426
rect 1052 350 1082 426
rect 1016 334 1082 350
rect 1016 300 1032 334
rect 1066 300 1082 334
rect 1016 284 1082 300
rect 1218 350 1248 426
rect 1218 334 1284 350
rect 1218 300 1234 334
rect 1268 300 1284 334
rect 1218 284 1284 300
rect 662 224 728 240
rect 878 234 974 250
rect 262 168 328 184
rect 262 134 278 168
rect 312 134 328 168
rect 262 118 328 134
rect 298 84 328 118
rect 464 168 530 184
rect 464 134 480 168
rect 514 134 530 168
rect 464 118 530 134
rect 572 168 638 184
rect 572 134 588 168
rect 622 134 638 168
rect 572 118 638 134
rect 464 84 494 118
rect 572 84 602 118
rect 680 84 710 224
rect 878 200 894 234
rect 928 200 974 234
rect 878 184 974 200
rect 1326 184 1356 426
rect 1434 350 1464 384
rect 1434 334 1500 350
rect 1434 300 1450 334
rect 1484 300 1500 334
rect 1434 284 1500 300
rect 944 84 974 184
rect 1016 168 1082 184
rect 1016 134 1032 168
rect 1066 134 1082 168
rect 1016 118 1082 134
rect 1052 84 1082 118
rect 1218 168 1284 184
rect 1218 134 1234 168
rect 1268 134 1284 168
rect 1218 118 1284 134
rect 1326 168 1392 184
rect 1326 134 1342 168
rect 1376 134 1392 168
rect 1326 118 1392 134
rect 1218 84 1248 118
rect 1326 84 1356 118
rect 1434 84 1464 284
rect 190 -30 220 0
rect 298 -30 328 0
rect 464 -30 494 0
rect 572 -30 602 0
rect 680 -30 710 0
rect 944 -30 974 0
rect 1052 -30 1082 0
rect 1218 -30 1248 0
rect 1326 -30 1356 0
rect 1434 -30 1464 0
rect 0 -72 30 -42
<< polycont >>
rect 278 300 312 334
rect 480 300 514 334
rect -50 216 -16 250
rect 170 202 204 236
rect 678 240 712 274
rect 1032 300 1066 334
rect 1234 300 1268 334
rect 278 134 312 168
rect 480 134 514 168
rect 588 134 622 168
rect 894 200 928 234
rect 1450 300 1484 334
rect 1032 134 1066 168
rect 1234 134 1268 168
rect 1342 134 1376 168
<< locali >>
rect -98 678 1612 697
rect -98 636 248 678
rect 282 636 448 678
rect 482 636 648 678
rect 682 636 848 678
rect 882 636 1048 678
rect 1082 636 1248 678
rect 1282 636 1448 678
rect 1482 636 1612 678
rect -45 536 -11 636
rect -45 384 -11 400
rect 41 536 75 552
rect 145 492 179 636
rect 145 426 179 458
rect 379 494 413 552
rect -66 250 0 266
rect -66 216 -50 250
rect -16 216 0 250
rect -66 200 0 216
rect 41 152 75 400
rect 262 334 328 350
rect 262 300 278 334
rect 312 300 328 334
rect 262 284 328 300
rect 379 257 413 460
rect 624 494 658 636
rect 624 384 658 460
rect 780 494 814 552
rect 464 334 530 350
rect 464 300 480 334
rect 514 300 530 334
rect 464 284 530 300
rect 662 274 728 290
rect 154 236 220 252
rect 154 202 170 236
rect 204 202 220 236
rect 154 186 220 202
rect 367 245 425 257
rect 367 211 379 245
rect 413 211 425 245
rect 662 240 678 274
rect 712 240 728 274
rect 662 224 728 240
rect 780 234 814 460
rect 899 494 933 636
rect 899 384 933 460
rect 1133 494 1167 552
rect 1016 334 1082 350
rect 1016 300 1032 334
rect 1066 300 1082 334
rect 1016 284 1082 300
rect 878 234 944 250
rect 367 199 425 211
rect 780 200 894 234
rect 928 200 944 234
rect 262 168 328 184
rect 262 152 278 168
rect 41 134 278 152
rect 312 134 328 168
rect 41 118 328 134
rect -45 68 -11 84
rect -45 -84 -11 16
rect 41 68 75 118
rect 41 0 75 16
rect 145 68 179 84
rect 145 -84 179 16
rect 379 68 413 199
rect 379 0 413 16
rect 464 168 530 184
rect 464 134 480 168
rect 514 134 530 168
rect 464 118 530 134
rect 572 168 638 184
rect 572 134 588 168
rect 622 152 638 168
rect 780 152 814 200
rect 878 184 944 200
rect 622 134 814 152
rect 572 118 814 134
rect 1016 168 1082 184
rect 1016 134 1032 168
rect 1066 134 1082 168
rect 1016 118 1082 134
rect 464 22 498 118
rect 624 68 658 84
rect 464 10 522 22
rect 464 -24 476 10
rect 510 -24 522 10
rect 464 -36 522 -24
rect 624 -84 658 16
rect 780 68 814 118
rect 780 0 814 16
rect 899 68 933 84
rect 899 -84 933 16
rect 1133 68 1167 460
rect 1378 494 1412 636
rect 1378 384 1412 460
rect 1534 494 1568 552
rect 1218 334 1284 350
rect 1218 300 1234 334
rect 1268 300 1284 334
rect 1218 284 1284 300
rect 1434 334 1500 350
rect 1434 300 1450 334
rect 1484 300 1500 334
rect 1434 284 1500 300
rect 1218 168 1284 184
rect 1218 134 1234 168
rect 1268 134 1284 168
rect 1218 118 1284 134
rect 1326 168 1392 184
rect 1326 134 1342 168
rect 1376 152 1392 168
rect 1534 152 1568 460
rect 1376 134 1568 152
rect 1326 118 1568 134
rect 1378 68 1412 84
rect 1167 46 1225 58
rect 1167 16 1179 46
rect 1133 12 1179 16
rect 1213 12 1225 46
rect 1133 0 1225 12
rect 1378 -84 1412 16
rect 1534 68 1568 118
rect 1534 0 1568 16
rect -98 -103 248 -84
rect -98 -145 48 -103
rect 82 -126 248 -103
rect 282 -126 448 -84
rect 482 -126 648 -84
rect 682 -126 848 -84
rect 882 -126 1048 -84
rect 1082 -126 1248 -84
rect 1282 -126 1448 -84
rect 1482 -126 1612 -84
rect 82 -145 1612 -126
<< viali >>
rect 248 670 282 678
rect 248 644 282 670
rect 448 670 482 678
rect 448 644 482 670
rect 648 670 682 678
rect 648 644 682 670
rect 848 670 882 678
rect 848 644 882 670
rect 1048 670 1082 678
rect 1048 644 1082 670
rect 1248 670 1282 678
rect 1248 644 1282 670
rect 1448 670 1482 678
rect 1448 644 1482 670
rect -50 216 -16 250
rect 278 300 312 334
rect 480 300 514 334
rect 170 202 204 236
rect 379 211 413 245
rect 678 240 712 274
rect 1032 300 1066 334
rect 278 134 312 168
rect 480 134 514 168
rect 1032 134 1066 168
rect 476 -24 510 10
rect 1234 300 1268 334
rect 1450 300 1484 334
rect 1234 134 1268 168
rect 1179 12 1213 46
rect 1534 16 1568 50
rect 48 -111 82 -103
rect 48 -137 82 -111
rect 248 -118 282 -92
rect 248 -126 282 -118
rect 448 -118 482 -92
rect 448 -126 482 -118
rect 648 -118 682 -92
rect 648 -126 682 -118
rect 848 -118 882 -92
rect 848 -126 882 -118
rect 1048 -118 1082 -92
rect 1048 -126 1082 -118
rect 1248 -118 1282 -92
rect 1248 -126 1282 -118
rect 1448 -118 1482 -92
rect 1448 -126 1482 -118
<< metal1 >>
rect -98 678 1612 697
rect -98 644 248 678
rect 282 644 448 678
rect 482 644 648 678
rect 682 644 848 678
rect 882 644 1048 678
rect 1082 644 1248 678
rect 1282 644 1448 678
rect 1482 644 1612 678
rect -98 636 1612 644
rect -50 384 1268 418
rect -50 262 -16 384
rect 278 346 312 384
rect 464 346 1066 350
rect 1234 346 1268 384
rect 266 334 324 346
rect 266 300 278 334
rect 312 300 324 334
rect 464 334 1078 346
rect 464 316 480 334
rect 266 288 324 300
rect 468 300 480 316
rect 514 316 1032 334
rect 514 300 526 316
rect 468 288 526 300
rect 1020 300 1032 316
rect 1066 316 1078 334
rect 1222 334 1280 346
rect 1066 308 1128 316
rect 1066 300 1134 308
rect 1020 288 1134 300
rect 1222 300 1234 334
rect 1268 300 1280 334
rect 1222 288 1280 300
rect 1438 334 1496 346
rect 1438 300 1450 334
rect 1484 300 1496 334
rect 1438 288 1496 300
rect 126 268 216 280
rect -94 250 -4 262
rect -94 184 -82 250
rect -16 184 -4 250
rect 126 202 138 268
rect 204 202 216 268
rect 666 274 724 286
rect 126 190 216 202
rect 367 245 425 257
rect 666 245 678 274
rect 367 211 379 245
rect 413 240 678 245
rect 712 240 724 274
rect 413 228 724 240
rect 413 211 711 228
rect 367 199 425 211
rect -94 172 -4 184
rect -50 22 -16 172
rect 266 168 324 180
rect 266 134 278 168
rect 312 134 324 168
rect 266 122 324 134
rect 468 168 526 180
rect 468 134 480 168
rect 514 152 526 168
rect 1020 168 1078 180
rect 1020 152 1032 168
rect 514 134 1032 152
rect 1066 134 1078 168
rect 468 122 1078 134
rect 1106 140 1134 288
rect 1222 168 1280 180
rect 1222 140 1234 168
rect 1106 134 1234 140
rect 1268 134 1280 168
rect 1106 122 1280 134
rect 278 84 312 122
rect 524 118 1064 122
rect 1106 106 1252 122
rect 1106 84 1134 106
rect 278 50 1134 84
rect 1167 56 1225 58
rect 1438 56 1466 288
rect 1528 72 1596 78
rect 1528 62 1534 72
rect 1167 46 1466 56
rect -50 10 522 22
rect -50 -12 476 10
rect 464 -24 476 -12
rect 510 -24 522 10
rect 1167 12 1179 46
rect 1213 22 1466 46
rect 1213 12 1225 22
rect 1167 0 1225 12
rect 1522 16 1534 62
rect 1590 16 1596 72
rect 1522 10 1596 16
rect 1522 4 1580 10
rect 464 -36 522 -24
rect -98 -92 1612 -84
rect -98 -103 248 -92
rect -98 -137 48 -103
rect 82 -126 248 -103
rect 282 -126 448 -92
rect 482 -126 648 -92
rect 682 -126 848 -92
rect 882 -126 1048 -92
rect 1082 -126 1248 -92
rect 1282 -126 1448 -92
rect 1482 -126 1612 -92
rect 82 -137 1612 -126
rect -98 -145 1612 -137
<< via1 >>
rect -82 216 -50 250
rect -50 216 -16 250
rect -82 184 -16 216
rect 138 236 204 268
rect 138 202 170 236
rect 170 202 204 236
rect 1534 50 1590 72
rect 1534 16 1568 50
rect 1568 16 1590 50
<< metal2 >>
rect 126 268 216 280
rect -94 250 -4 262
rect -94 184 -82 250
rect -16 184 -4 250
rect 126 202 138 268
rect 204 202 216 268
rect 126 190 216 202
rect -94 172 -4 184
rect 1528 72 1596 78
rect 1528 16 1534 72
rect 1590 16 1596 72
rect 1528 10 1596 16
<< labels >>
rlabel metal2 170 202 204 236 5 D
port 2 s
rlabel metal2 1534 16 1590 72 5 Q
port 3 s
rlabel locali -68 -119 -68 -119 5 gnd
rlabel locali -50 670 -50 670 5 vdd
rlabel locali 58 136 58 136 5 CLK_n
rlabel viali 396 228 396 228 5 common_1
rlabel locali 800 218 800 218 5 inverter_1_out
rlabel viali 1196 30 1196 30 5 common_2
rlabel metal2 -50 216 -16 250 5 CLK
port 1 s
<< end >>
