* NGSPICE file created from buffer_fo4.ext - technology: sky130A

.subckt buffer_fo4 A B gnd vdd
X0 a_n240_0# A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
X1 B a_n240_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.47 pd=3.92 as=0.504 ps=3.96 w=1.68 l=0.15
X2 a_n240_0# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X3 vdd a_n240_0# B vdd sky130_fd_pr__pfet_01v8 ad=1.01 pd=7.32 as=0.941 ps=7.28 w=3.36 l=0.15
.ends

