* NGSPICE file created from register.ext - technology: sky130A

.subckt d_flip_flop CLK D Q gnd vdd a_494_0# a_1248_0# CLK_n a_220_0# inverter_1_out
+ common_2 common_1 a_974_0#
X0 inverter_1_out common_1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X1 gnd inverter_1_out a_494_0# gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
X2 common_2 CLK_n a_974_426# vdd sky130_fd_pr__pfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 gnd Q a_1248_0# gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
X4 a_974_0# inverter_1_out gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X5 a_220_426# D vdd vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X6 a_494_0# CLK common_1 gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X7 a_1248_0# CLK_n common_2 gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X8 CLK_n CLK vdd vdd sky130_fd_pr__pfet_01v8 ad=0.445 pd=3.89 as=0.445 ps=3.89 w=1.68 l=0.15
X9 common_1 CLK a_220_426# vdd sky130_fd_pr__pfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X10 Q common_2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.34 pd=2.8 as=0.134 ps=1.23 w=0.84 l=0.15
X11 a_1248_426# CLK common_2 vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X12 CLK_n CLK gnd gnd sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
X13 common_1 CLK_n a_220_0# gnd sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X14 vdd Q a_1248_426# vdd sky130_fd_pr__pfet_01v8 ad=0.134 pd=1.23 as=0.0819 ps=0.81 w=0.42 l=0.15
X15 common_2 CLK a_974_0# gnd sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X16 inverter_1_out common_1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X17 Q common_2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X18 a_494_426# CLK_n common_1 vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X19 a_974_426# inverter_1_out vdd vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X20 a_220_0# D gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X21 vdd inverter_1_out a_494_426# vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
C0 inverter_1_out common_2 0.0217f
C1 CLK_n vdd 0.318f
C2 common_1 CLK_n 0.257f
C3 Q vdd 0.172f
C4 Q common_1 2.17e-19
C5 a_220_426# vdd 0.00638f
C6 inverter_1_out CLK_n 0.21f
C7 a_220_426# common_1 0.00211f
C8 a_494_426# CLK_n 0.00166f
C9 inverter_1_out Q 0.00505f
C10 common_1 vdd 0.175f
C11 CLK D 0.188f
C12 inverter_1_out vdd 0.302f
C13 inverter_1_out common_1 0.241f
C14 a_494_426# vdd 0.00747f
C15 a_1248_426# CLK 0.0028f
C16 a_494_426# common_1 0.00211f
C17 CLK common_2 0.116f
C18 a_220_0# common_2 9.78e-20
C19 CLK CLK_n 1.39f
C20 a_220_0# CLK_n 0.00636f
C21 CLK Q 0.0622f
C22 a_220_0# Q 1.24e-19
C23 CLK a_220_426# 0.00458f
C24 CLK vdd 0.661f
C25 CLK common_1 0.294f
C26 a_220_0# common_1 0.00135f
C27 CLK inverter_1_out 0.224f
C28 CLK a_494_426# 0.00292f
C29 common_2 a_494_0# 2.69e-19
C30 common_2 a_974_0# 0.00277f
C31 CLK_n a_494_0# 0.00356f
C32 Q a_494_0# 1.34e-19
C33 CLK_n a_974_0# 0.00401f
C34 a_974_426# common_2 0.00211f
C35 vdd a_494_0# 2.34e-19
C36 Q a_974_0# 3.81e-19
C37 a_220_0# CLK 0.00497f
C38 common_2 a_1248_0# 0.00945f
C39 vdd a_974_0# 2.34e-19
C40 a_974_426# CLK_n 0.00166f
C41 CLK_n a_1248_0# 0.00313f
C42 Q a_1248_0# 9.54e-19
C43 a_974_426# vdd 0.00744f
C44 common_2 D 1.9e-19
C45 a_1248_426# common_2 0.00273f
C46 vdd a_1248_0# 3.63e-19
C47 D CLK_n 0.122f
C48 Q D 2.13e-19
C49 CLK a_494_0# 0.00903f
C50 common_2 CLK_n 0.209f
C51 D vdd 0.109f
C52 D common_1 0.0338f
C53 common_2 Q 0.269f
C54 CLK a_974_0# 0.00228f
C55 a_1248_426# vdd 0.00627f
C56 inverter_1_out D 0.00602f
C57 common_2 vdd 0.165f
C58 common_2 common_1 3.81e-19
C59 Q CLK_n 0.0719f
C60 CLK a_974_426# 0.00292f
C61 a_220_426# CLK_n 6.84e-19
C62 Q gnd 0.492f
C63 D gnd 0.27f
C64 CLK gnd 1.15f
C65 vdd gnd 2.63f
C66 a_1248_0# gnd 0.00421f
C67 a_974_0# gnd 0.00647f
C68 a_494_0# gnd 0.00449f
C69 a_220_0# gnd 0.00356f
C70 a_1248_426# gnd 2.68e-19
C71 a_974_426# gnd 2.68e-19
C72 a_494_426# gnd 2.68e-19
C73 common_2 gnd 0.517f
C74 common_1 gnd 0.302f
C75 inverter_1_out gnd 0.593f
C76 CLK_n gnd 0.855f
.ends

.subckt and2 A B Y gnd vdd a_30_n42# Y_n
X0 vdd B Y_n vdd sky130_fd_pr__pfet_01v8 ad=0.212 pd=1.35 as=0.118 ps=1.12 w=0.84 l=0.15
X1 Y Y_n vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.212 ps=1.35 w=0.84 l=0.15
X2 Y Y_n gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.159 ps=1.35 w=0.42 l=0.15
X3 Y_n A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X4 gnd B a_30_n42# gnd sky130_fd_pr__nfet_01v8 ad=0.159 pd=1.35 as=0.118 ps=1.12 w=0.84 l=0.15
X5 a_30_n42# A Y_n gnd sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
C0 Y_n vdd 0.186f
C1 A Y 0.00134f
C2 B Y 0.0233f
C3 A B 0.0938f
C4 a_30_n42# Y 9.31e-19
C5 Y_n Y 0.0794f
C6 A Y_n 0.0914f
C7 vdd Y 0.0836f
C8 A vdd 0.072f
C9 Y_n B 0.176f
C10 vdd B 0.108f
C11 Y_n a_30_n42# 0.0116f
C12 a_30_n42# vdd 4.51e-19
C13 Y gnd 0.284f
C14 B gnd 0.248f
C15 A gnd 0.322f
C16 vdd gnd 0.757f
C17 a_30_n42# gnd 0.00713f
C18 Y_n gnd 0.444f
.ends

.subckt register D CLK EN Q gnd vdd
Xd_flip_flop_0 and2_0/Y D Q gnd vdd d_flip_flop_0/a_494_0# d_flip_flop_0/a_1248_0#
+ d_flip_flop_0/CLK_n d_flip_flop_0/a_220_0# d_flip_flop_0/inverter_1_out d_flip_flop_0/common_2
+ d_flip_flop_0/common_1 d_flip_flop_0/a_974_0# d_flip_flop
Xand2_0 CLK EN and2_0/Y gnd vdd and2_0/a_30_n42# and2_0/Y_n and2
C0 CLK and2_0/Y 0.0199f
C1 d_flip_flop_0/inverter_1_out EN 1.44e-19
C2 and2_0/a_30_n42# and2_0/Y 7.24e-19
C3 EN Q 2.99e-20
C4 and2_0/Y_n D 0.00817f
C5 D EN 7.78e-19
C6 vdd D 0.00388f
C7 d_flip_flop_0/CLK_n and2_0/Y 0.0351f
C8 CLK D 4.88e-20
C9 d_flip_flop_0/common_2 EN 3.89e-20
C10 vdd and2_0/Y_n 0.014f
C11 vdd EN 0.00216f
C12 and2_0/Y_n CLK 2.84e-32
C13 CLK EN -1.42e-32
C14 and2_0/Y d_flip_flop_0/a_220_0# 6.81e-19
C15 and2_0/Y d_flip_flop_0/a_494_0# 2.46e-19
C16 d_flip_flop_0/CLK_n and2_0/Y_n 5.91e-19
C17 d_flip_flop_0/a_1248_0# and2_0/Y 8.55e-20
C18 d_flip_flop_0/CLK_n EN 0.00102f
C19 d_flip_flop_0/CLK_n vdd 5.37e-19
C20 Q d_flip_flop_0/a_220_0# -1.39e-35
C21 d_flip_flop_0/common_1 and2_0/Y 9.82e-19
C22 and2_0/Y d_flip_flop_0/a_974_0# 1.25e-19
C23 d_flip_flop_0/inverter_1_out and2_0/Y 7.03e-19
C24 and2_0/Y Q 1.66e-19
C25 D and2_0/Y 0.00132f
C26 d_flip_flop_0/common_1 EN 2.23e-19
C27 d_flip_flop_0/common_2 and2_0/Y 3.33e-19
C28 and2_0/Y_n and2_0/Y 0.0383f
C29 and2_0/Y EN 0.0186f
C30 vdd and2_0/Y 0.0522f
C31 vdd gnd 3.28f
C32 EN gnd 0.231f
C33 CLK gnd 0.306f
C34 and2_0/a_30_n42# gnd 0.00713f
C35 and2_0/Y_n gnd 0.445f
C36 Q gnd 0.492f
C37 D gnd 0.257f
C38 and2_0/Y gnd 1.29f
C39 d_flip_flop_0/a_1248_0# gnd 0.00421f
C40 d_flip_flop_0/a_974_0# gnd 0.00647f
C41 d_flip_flop_0/a_494_0# gnd 0.00449f
C42 d_flip_flop_0/a_220_0# gnd 0.00356f
C43 d_flip_flop_0/a_1248_426# gnd 2.68e-19 $ **FLOATING
C44 d_flip_flop_0/a_974_426# gnd 2.68e-19 $ **FLOATING
C45 d_flip_flop_0/a_494_426# gnd 2.68e-19 $ **FLOATING
C46 d_flip_flop_0/common_2 gnd 0.517f
C47 d_flip_flop_0/common_1 gnd 0.302f
C48 d_flip_flop_0/inverter_1_out gnd 0.593f
C49 d_flip_flop_0/CLK_n gnd 0.855f
.ends

