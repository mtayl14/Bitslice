** sch_path: /home/mtayl14/Projects/Bitslice/xschem/mux21.sch
.subckt mux21 S A B Y
*.PININFO S:I A:I B:I Y:O
x1 S A Y net1 t_gate
x2 net1 B Y S t_gate
x3 net1 S inv
.ends

* expanding   symbol:  t_gate.sym # of pins=4
** sym_path: /home/mtayl14/Projects/Bitslice/xschem/t_gate.sym
** sch_path: /home/mtayl14/Projects/Bitslice/xschem/t_gate.sch
.subckt t_gate E_n in out E
*.PININFO in:I out:O E:I E_n:I
XM1 in E out GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 in E_n out VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  inv.sym # of pins=2
** sym_path: /home/mtayl14/Projects/Bitslice/xschem/inv.sym
** sch_path: /home/mtayl14/Projects/Bitslice/xschem/inv.sch
.subckt inv Z A
*.PININFO A:I Z:O
XM1 Z A GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Z A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.84 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
