../magic/datapath.spice