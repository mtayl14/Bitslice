magic
tech sky130A
magscale 1 2
timestamp 1701898898
<< locali >>
rect 541 681 575 697
rect 1841 534 1893 586
<< viali >>
rect 541 697 575 731
<< metal1 >>
rect 0 781 123 842
rect 332 736 398 742
rect 332 724 338 736
rect 52 690 338 724
rect 52 626 86 690
rect 332 682 338 690
rect 392 682 398 736
rect 529 731 802 749
rect 529 697 541 731
rect 575 721 802 731
rect 575 697 587 721
rect 529 685 587 697
rect 332 676 398 682
rect 23 620 89 626
rect 23 566 29 620
rect 83 566 89 620
rect 23 560 89 566
rect 774 488 802 721
rect 3416 694 3480 700
rect 3416 690 3422 694
rect 1842 654 3422 690
rect 1844 592 1878 654
rect 3416 642 3422 654
rect 3474 642 3480 694
rect 3416 636 3480 642
rect 1835 586 1899 592
rect 1835 534 1841 586
rect 1893 534 1899 586
rect 1835 528 1899 534
rect 2007 493 2071 499
rect 242 479 306 485
rect 242 427 248 479
rect 300 427 306 479
rect 2007 441 2013 493
rect 2065 441 2071 493
rect 2007 435 2071 441
rect 46 288 80 422
rect 242 421 306 427
rect 922 419 986 425
rect 922 367 928 419
rect 980 367 986 419
rect 2874 370 3170 398
rect 922 361 986 367
rect 772 345 836 351
rect 772 293 778 345
rect 830 293 836 345
rect 46 260 460 288
rect 772 287 836 293
rect 432 212 460 260
rect 142 162 166 164
rect 142 117 174 162
rect 628 117 658 162
rect 142 89 658 117
rect 0 0 121 61
<< via1 >>
rect 338 682 392 736
rect 29 566 83 620
rect 3422 642 3474 694
rect 1841 534 1893 586
rect 248 427 300 479
rect 2013 441 2065 493
rect 928 367 980 419
rect 778 293 830 345
<< metal2 >>
rect 23 620 89 626
rect 23 566 29 620
rect 83 566 89 620
rect 23 560 89 566
rect 248 485 300 930
rect 348 756 808 758
rect 348 742 810 756
rect 332 736 810 742
rect 332 682 338 736
rect 392 720 810 736
rect 392 682 398 720
rect 332 676 398 682
rect 242 479 306 485
rect 30 427 82 479
rect 242 427 248 479
rect 300 427 306 479
rect 242 421 306 427
rect 248 -70 300 421
rect 778 351 810 720
rect 924 682 976 930
rect 924 630 1696 682
rect 922 419 986 425
rect 922 367 928 419
rect 980 367 986 419
rect 922 361 986 367
rect 772 345 836 351
rect 772 293 778 345
rect 830 293 836 345
rect 772 287 836 293
rect 924 -70 976 361
rect 1644 310 1696 630
rect 1835 586 1899 592
rect 1835 534 1841 586
rect 1893 534 1899 586
rect 1835 528 1899 534
rect 2007 493 2071 499
rect 2007 441 2013 493
rect 2065 441 2071 493
rect 2007 435 2071 441
rect 2008 310 2060 435
rect 1644 258 2060 310
rect 2115 -70 2167 930
rect 3305 -70 3357 930
rect 3416 694 3480 700
rect 3416 642 3422 694
rect 3474 692 3480 694
rect 3474 654 3802 692
rect 3474 642 3480 654
rect 3416 636 3480 642
rect 3748 380 3802 654
rect 5146 161 5202 217
use addf  addf_0
timestamp 1701894535
transform 1 0 698 0 1 -20
box -18 0 1411 897
use buffer_fo4  buffer_fo4_0
timestamp 1701892857
transform 1 0 2453 0 1 145
box -368 -145 655 706
use inverter  inverter_0
timestamp 1701892814
transform 1 0 98 0 1 145
box -98 -145 128 706
use mux21  mux21_0
timestamp 1701892517
transform 1 0 310 0 1 145
box -100 -145 396 706
use register  register_0
timestamp 1701889381
transform 1 0 3080 0 1 0
box 0 0 2144 851
<< labels >>
rlabel metal1 0 0 121 61 5 gnd
port 0 s
rlabel metal1 0 781 123 842 5 vdd
port 1 s
rlabel metal2 30 427 82 479 5 B
port 3 s
rlabel via1 248 427 300 479 5 SUB
port 5 s
rlabel via1 778 293 830 345 5 A
port 4 s
rlabel metal2 928 367 980 419 5 CI
port 6 s
rlabel metal2 2013 441 2065 493 5 CO
port 9 s
rlabel metal2 2115 427 2167 479 5 CLK
port 8 s
rlabel metal2 3305 427 3357 479 5 STORE
port 7 s
rlabel metal2 5146 161 5202 217 5 Q
port 10 s
<< end >>
