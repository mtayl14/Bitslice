magic
tech sky130A
magscale 1 2
timestamp 1701892857
<< nwell >>
rect -368 342 655 706
<< nmos >>
rect -270 0 -240 84
rect 115 45 451 75
<< pmos >>
rect -270 384 -240 552
rect -53 434 619 464
<< ndiff >>
rect 115 120 451 131
rect -323 68 -270 84
rect -323 16 -315 68
rect -281 16 -270 68
rect -323 0 -270 16
rect -240 68 -187 84
rect -240 16 -229 68
rect -195 16 -187 68
rect 115 86 131 120
rect 435 86 451 120
rect 115 75 451 86
rect -240 0 -187 16
rect 115 30 451 45
rect 115 -4 131 30
rect 435 -4 451 30
rect 115 -15 451 -4
<< pdiff >>
rect -323 536 -270 552
rect -323 400 -315 536
rect -281 400 -270 536
rect -323 384 -270 400
rect -240 536 -187 552
rect -240 400 -229 536
rect -195 400 -187 536
rect -53 516 619 524
rect -53 475 -37 516
rect 603 475 619 516
rect -53 464 619 475
rect -240 384 -187 400
rect -53 423 619 434
rect -53 386 71 423
rect 603 386 619 423
rect -53 378 619 386
<< ndiffc >>
rect -315 16 -281 68
rect -229 16 -195 68
rect 131 86 435 120
rect 131 -4 435 30
<< pdiffc >>
rect -315 400 -281 536
rect -229 400 -195 536
rect -37 475 603 516
rect 71 386 603 423
<< psubdiff >>
rect -272 -118 -247 -84
rect -213 -118 -188 -84
rect -2 -118 23 -84
rect 57 -118 82 -84
rect 136 -118 161 -84
rect 195 -118 220 -84
rect 274 -118 299 -84
rect 333 -118 358 -84
rect 412 -118 437 -84
rect 471 -118 496 -84
<< nsubdiff >>
rect -270 636 -245 670
rect -211 636 -186 670
rect 0 636 25 670
rect 59 636 84 670
rect 138 636 163 670
rect 197 636 222 670
rect 276 636 301 670
rect 335 636 360 670
rect 414 636 439 670
rect 473 636 498 670
<< psubdiffcont >>
rect -247 -118 -213 -84
rect 23 -118 57 -84
rect 161 -118 195 -84
rect 299 -118 333 -84
rect 437 -118 471 -84
<< nsubdiffcont >>
rect -245 636 -211 670
rect 25 636 59 670
rect 163 636 197 670
rect 301 636 335 670
rect 439 636 473 670
<< poly >>
rect -270 552 -240 582
rect -153 448 -53 464
rect -153 414 -137 448
rect -103 434 -53 448
rect 619 434 649 464
rect -103 414 -87 434
rect -153 398 -87 414
rect -270 350 -240 384
rect -336 334 -240 350
rect -336 300 -320 334
rect -286 300 -240 334
rect -336 284 -240 300
rect -270 84 -240 284
rect 15 95 81 111
rect 15 61 31 95
rect 65 75 81 95
rect 65 61 115 75
rect 15 45 115 61
rect 451 45 481 75
rect -270 -30 -240 0
<< polycont >>
rect -137 414 -103 448
rect -320 300 -286 334
rect 31 61 65 95
<< locali >>
rect -368 678 655 697
rect -368 636 -245 678
rect -211 636 25 678
rect 59 636 163 678
rect 197 636 301 678
rect 335 636 439 678
rect 473 636 655 678
rect -315 536 -281 636
rect -315 384 -281 400
rect -229 536 -195 552
rect -53 516 619 636
rect -53 475 -37 516
rect 603 475 619 516
rect -53 468 619 475
rect -195 448 -87 464
rect -195 414 -137 448
rect -103 414 -87 448
rect -195 400 -87 414
rect -336 334 -270 350
rect -336 300 -320 334
rect -286 300 -270 334
rect -336 284 -270 300
rect -229 92 -87 400
rect 55 423 619 434
rect 55 386 71 423
rect 603 386 619 423
rect 55 378 619 386
rect 115 262 451 378
rect 115 228 398 262
rect 432 228 451 262
rect 115 120 451 228
rect 15 95 81 111
rect 15 92 31 95
rect -315 68 -281 84
rect -315 -84 -281 16
rect -229 68 31 92
rect -195 61 31 68
rect 65 61 81 95
rect 115 86 131 120
rect 435 86 451 120
rect 115 75 451 86
rect -195 58 81 61
rect 15 45 81 58
rect -229 0 -195 16
rect 115 30 451 41
rect 115 -4 131 30
rect 435 -4 451 30
rect 115 -84 451 -4
rect -368 -126 -247 -84
rect -213 -126 23 -84
rect 57 -126 161 -84
rect 195 -126 299 -84
rect 333 -126 437 -84
rect 471 -126 653 -84
rect -368 -145 653 -126
<< viali >>
rect -245 670 -211 678
rect -245 644 -211 670
rect 25 670 59 678
rect 25 644 59 670
rect 163 670 197 678
rect 163 644 197 670
rect 301 670 335 678
rect 301 644 335 670
rect 439 670 473 678
rect 439 644 473 670
rect -320 300 -286 334
rect 398 228 432 262
rect -247 -118 -213 -92
rect -247 -126 -213 -118
rect 23 -118 57 -92
rect 23 -126 57 -118
rect 161 -118 195 -92
rect 161 -126 195 -118
rect 299 -118 333 -92
rect 299 -126 333 -118
rect 437 -118 471 -92
rect 437 -126 471 -118
<< metal1 >>
rect -368 678 655 697
rect -368 644 -245 678
rect -211 644 25 678
rect 59 644 163 678
rect 197 644 301 678
rect 335 644 439 678
rect 473 644 655 678
rect -368 636 655 644
rect -332 340 -274 346
rect -344 334 -274 340
rect -344 282 -338 334
rect -286 288 -274 334
rect -286 282 -280 288
rect -344 276 -280 282
rect 383 271 447 277
rect 383 219 389 271
rect 441 219 447 271
rect 383 213 447 219
rect -368 -92 653 -84
rect -368 -126 -247 -92
rect -213 -126 23 -92
rect 57 -126 161 -92
rect 195 -126 299 -92
rect 333 -126 437 -92
rect 471 -126 653 -92
rect -368 -145 653 -126
<< via1 >>
rect -338 300 -320 334
rect -320 300 -286 334
rect -338 282 -286 300
rect 389 262 441 271
rect 389 228 398 262
rect 398 228 432 262
rect 432 228 441 262
rect 389 219 441 228
<< metal2 >>
rect -344 334 -280 340
rect -344 282 -338 334
rect -286 282 -280 334
rect -344 276 -280 282
rect 383 271 447 277
rect 383 219 389 271
rect 441 219 447 271
rect 383 213 447 219
<< labels >>
rlabel via1 416 246 416 246 5 B
port 2 s
rlabel metal1 -124 -110 -124 -110 5 gnd
rlabel metal1 -128 666 -128 666 5 vdd
rlabel via1 -312 308 -312 308 5 A
port 1 s
rlabel metal1 -348 664 -348 664 5 vdd
port 4 s
rlabel metal1 -346 -116 -346 -116 5 gnd
port 3 s
<< end >>
