magic
tech sky130A
magscale 1 2
timestamp 1701892517
<< nwell >>
rect -98 348 396 706
<< nmos >>
rect 0 0 30 84
rect 190 0 220 84
rect 276 0 306 84
<< pmos >>
rect 0 384 30 552
rect 190 384 220 552
rect 276 384 306 552
<< ndiff >>
rect -53 68 0 84
rect -53 16 -45 68
rect -11 16 0 68
rect -53 0 0 16
rect 30 68 83 84
rect 30 16 41 68
rect 75 16 83 68
rect 30 0 83 16
rect 137 68 190 84
rect 137 16 145 68
rect 179 16 190 68
rect 137 0 190 16
rect 220 68 276 84
rect 220 16 231 68
rect 265 16 276 68
rect 220 0 276 16
rect 306 68 359 84
rect 306 16 317 68
rect 351 16 359 68
rect 306 0 359 16
<< pdiff >>
rect -53 536 0 552
rect -53 400 -45 536
rect -11 400 0 536
rect -53 384 0 400
rect 30 536 83 552
rect 30 400 41 536
rect 75 400 83 536
rect 30 384 83 400
rect 137 536 190 552
rect 137 400 145 536
rect 179 400 190 536
rect 137 384 190 400
rect 220 536 276 552
rect 220 400 231 536
rect 265 400 276 536
rect 220 384 276 400
rect 306 536 359 552
rect 306 400 317 536
rect 351 400 359 536
rect 306 384 359 400
<< ndiffc >>
rect -45 16 -11 68
rect 41 16 75 68
rect 145 16 179 68
rect 231 16 265 68
rect 317 16 351 68
<< pdiffc >>
rect -45 400 -11 536
rect 41 400 75 536
rect 145 400 179 536
rect 231 400 265 536
rect 317 400 351 536
<< psubdiff >>
rect -2 -118 23 -84
rect 57 -118 82 -84
rect 136 -118 161 -84
rect 195 -118 220 -84
rect 274 -118 299 -84
rect 333 -118 358 -84
<< nsubdiff >>
rect 0 636 25 670
rect 59 636 84 670
rect 138 636 163 670
rect 197 636 222 670
rect 276 636 301 670
rect 335 636 360 670
<< psubdiffcont >>
rect 23 -118 57 -84
rect 161 -118 195 -84
rect 299 -118 333 -84
<< nsubdiffcont >>
rect 25 636 59 670
rect 163 636 197 670
rect 301 636 335 670
<< poly >>
rect 0 552 30 582
rect 190 552 220 582
rect 276 552 306 582
rect 0 350 30 384
rect 190 350 220 384
rect -60 334 30 350
rect -60 300 -44 334
rect -10 300 30 334
rect -60 284 30 300
rect 131 334 220 350
rect 131 300 147 334
rect 181 300 220 334
rect 131 284 220 300
rect 276 350 306 384
rect 276 334 365 350
rect 276 300 315 334
rect 349 300 365 334
rect 276 284 365 300
rect 0 84 30 284
rect 131 174 220 190
rect 131 140 147 174
rect 181 140 220 174
rect 131 124 220 140
rect 190 84 220 124
rect 276 174 365 190
rect 276 140 315 174
rect 349 140 365 174
rect 276 124 365 140
rect 276 84 306 124
rect 0 -30 30 0
rect 190 -30 220 0
rect 276 -30 306 0
<< polycont >>
rect -44 300 -10 334
rect 147 300 181 334
rect 315 300 349 334
rect 147 140 181 174
rect 315 140 349 174
<< locali >>
rect -98 678 396 697
rect -98 636 25 678
rect 59 636 163 678
rect 197 636 301 678
rect 335 636 396 678
rect -45 536 -11 636
rect -45 384 -11 400
rect 41 536 75 552
rect -60 334 6 350
rect -60 300 -44 334
rect -10 300 6 334
rect -60 284 6 300
rect 41 158 75 400
rect 145 536 179 552
rect 145 384 179 400
rect 231 536 265 552
rect 131 334 197 350
rect 131 300 147 334
rect 181 300 197 334
rect 131 284 197 300
rect 131 174 197 190
rect 131 158 147 174
rect 41 140 147 158
rect 181 140 197 174
rect 41 124 197 140
rect -45 68 -11 84
rect -45 -84 -11 16
rect 41 68 75 124
rect 41 0 75 16
rect 145 68 179 84
rect 145 0 179 16
rect 231 68 265 400
rect 317 536 351 552
rect 317 384 351 400
rect 299 334 365 350
rect 299 300 315 334
rect 349 300 365 334
rect 299 284 365 300
rect 299 174 365 190
rect 299 140 315 174
rect 349 140 365 174
rect 299 124 365 140
rect 231 0 265 16
rect 317 68 351 84
rect 317 0 351 16
rect -100 -126 23 -84
rect 57 -126 161 -84
rect 195 -126 299 -84
rect 333 -126 394 -84
rect -100 -145 394 -126
<< viali >>
rect 25 670 59 678
rect 25 644 59 670
rect 163 670 197 678
rect 163 644 197 670
rect 301 670 335 678
rect 301 644 335 670
rect 41 400 75 434
rect -44 300 -10 334
rect 145 502 179 536
rect 147 300 181 334
rect 41 34 75 68
rect 145 16 179 68
rect 317 502 351 536
rect 315 300 349 334
rect 315 140 349 174
rect 231 16 265 68
rect 317 16 351 68
rect 23 -118 57 -92
rect 23 -126 57 -118
rect 161 -118 195 -92
rect 161 -126 195 -118
rect 299 -118 333 -92
rect 299 -126 333 -118
<< metal1 >>
rect -98 678 396 697
rect -98 644 25 678
rect 59 644 163 678
rect 197 644 301 678
rect 335 644 396 678
rect -98 636 396 644
rect 133 542 191 548
rect 121 536 191 542
rect 121 484 127 536
rect 179 490 191 536
rect 305 542 363 548
rect 305 536 375 542
rect 305 490 317 536
rect 179 484 185 490
rect 121 478 185 484
rect 311 484 317 490
rect 369 484 375 536
rect 311 478 375 484
rect 29 440 87 446
rect 29 434 330 440
rect 29 400 41 434
rect 75 410 330 434
rect 75 400 87 410
rect 29 388 87 400
rect 300 350 330 410
rect 300 346 360 350
rect -56 340 2 346
rect 135 340 193 346
rect 300 340 361 346
rect -56 334 193 340
rect -56 300 -44 334
rect -10 310 147 334
rect -10 300 2 310
rect -56 288 2 300
rect 135 300 147 310
rect 181 300 193 334
rect 135 288 193 300
rect 303 334 361 340
rect 303 300 315 334
rect 349 300 361 334
rect 303 288 361 300
rect 163 250 193 288
rect 163 220 340 250
rect 310 186 340 220
rect 303 174 361 186
rect 303 140 315 174
rect 349 140 361 174
rect 303 128 361 140
rect 29 68 87 80
rect 133 74 191 80
rect 29 34 41 68
rect 75 34 87 68
rect 29 22 87 34
rect 121 68 191 74
rect 121 16 127 68
rect 179 16 191 68
rect 121 10 191 16
rect 133 4 191 10
rect 219 68 277 80
rect 219 16 222 68
rect 274 16 277 68
rect 219 4 277 16
rect 305 74 363 80
rect 305 68 375 74
rect 305 16 317 68
rect 369 16 375 68
rect 305 10 375 16
rect 305 4 363 10
rect -100 -92 394 -84
rect -100 -126 23 -92
rect 57 -126 161 -92
rect 195 -126 299 -92
rect 333 -126 394 -92
rect -100 -145 394 -126
<< via1 >>
rect 127 502 145 536
rect 145 502 179 536
rect 127 484 179 502
rect 317 502 351 536
rect 351 502 369 536
rect 317 484 369 502
rect 127 16 145 68
rect 145 16 179 68
rect 222 16 231 68
rect 231 16 265 68
rect 265 16 274 68
rect 317 16 351 68
rect 351 16 369 68
<< metal2 >>
rect 121 536 185 542
rect 121 484 127 536
rect 179 484 185 536
rect 121 478 185 484
rect 311 536 375 542
rect 311 484 317 536
rect 369 484 375 536
rect 311 478 375 484
rect 130 74 170 478
rect 330 74 370 478
rect 121 68 185 74
rect 121 16 127 68
rect 179 16 185 68
rect 121 10 185 16
rect 216 68 280 74
rect 216 16 222 68
rect 274 16 280 68
rect 216 10 280 16
rect 311 68 375 74
rect 311 16 317 68
rect 369 16 375 68
rect 311 10 375 16
<< labels >>
rlabel via1 248 42 248 42 5 Y
port 3 s
rlabel locali 60 140 60 140 5 S_n
rlabel via1 162 42 162 42 5 A
port 1 s
rlabel via1 334 42 334 42 5 B
port 2 s
rlabel viali 40 -101 40 -101 5 gnd
port 5 s
rlabel viali 42 653 42 653 1 vdd
port 6 n
rlabel viali -27 317 -27 317 5 S
port 4 s
rlabel viali 180 653 180 653 1 vdd
rlabel viali 318 653 318 653 1 vdd
rlabel viali 178 -101 178 -101 5 gnd
rlabel viali 316 -101 316 -101 5 gnd
<< end >>
