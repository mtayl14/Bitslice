magic
tech sky130A
magscale 1 2
timestamp 1701820176
<< nwell >>
rect -98 348 128 706
<< nmos >>
rect 0 0 30 84
<< pmos >>
rect 0 384 30 552
<< ndiff >>
rect -53 68 0 84
rect -53 16 -45 68
rect -11 16 0 68
rect -53 0 0 16
rect 30 68 83 84
rect 30 16 41 68
rect 75 16 83 68
rect 30 0 83 16
<< pdiff >>
rect -53 536 0 552
rect -53 400 -45 536
rect -11 400 0 536
rect -53 384 0 400
rect 30 536 83 552
rect 30 400 41 536
rect 75 400 83 536
rect 30 384 83 400
<< ndiffc >>
rect -45 16 -11 68
rect 41 16 75 68
<< pdiffc >>
rect -45 400 -11 536
rect 41 400 75 536
<< psubdiff >>
rect -2 -118 23 -84
rect 57 -118 82 -84
<< nsubdiff >>
rect 0 636 25 670
rect 59 636 84 670
<< psubdiffcont >>
rect 23 -118 57 -84
<< nsubdiffcont >>
rect 25 636 59 670
<< poly >>
rect 0 552 30 582
rect 0 350 30 384
rect -66 334 30 350
rect -66 300 -50 334
rect -16 300 30 334
rect -66 284 30 300
rect 0 84 30 284
rect 0 -30 30 0
<< polycont >>
rect -50 300 -16 334
<< locali >>
rect -98 678 128 697
rect -98 636 25 678
rect 59 636 128 678
rect -45 536 -11 636
rect -45 384 -11 400
rect 41 536 75 552
rect -66 334 0 350
rect -66 300 -50 334
rect -16 300 0 334
rect -66 284 0 300
rect -45 68 -11 84
rect 41 80 75 400
rect -45 -84 -11 16
rect 29 68 87 80
rect 29 16 41 68
rect 75 16 87 68
rect 29 4 87 16
rect 41 0 75 4
rect -98 -126 23 -84
rect 57 -126 126 -84
rect -98 -145 126 -126
<< viali >>
rect 25 670 59 678
rect 25 644 59 670
rect -50 300 -16 334
rect 41 16 75 68
rect 23 -118 57 -92
rect 23 -126 57 -118
<< metal1 >>
rect -98 678 128 697
rect -98 644 25 678
rect 59 644 128 678
rect -98 636 128 644
rect -62 340 -4 346
rect -74 334 -4 340
rect -74 282 -68 334
rect -16 288 -4 334
rect -16 282 -10 288
rect -74 276 -10 282
rect 29 74 87 80
rect 29 68 99 74
rect 29 16 41 68
rect 93 16 99 68
rect 29 10 99 16
rect 29 4 87 10
rect -98 -92 126 -84
rect -98 -126 23 -92
rect 57 -126 126 -92
rect -98 -145 126 -126
<< via1 >>
rect -68 300 -50 334
rect -50 300 -16 334
rect -68 282 -16 300
rect 41 16 75 68
rect 75 16 93 68
<< metal2 >>
rect -74 334 -10 340
rect -74 282 -68 334
rect -16 282 -10 334
rect -74 276 -10 282
rect 35 68 99 74
rect 35 16 41 68
rect 93 16 99 68
rect 35 10 99 16
<< labels >>
rlabel via1 -42 308 -42 308 5 A
port 1 s
rlabel via1 67 42 67 42 5 B
port 2 s
rlabel metal1 -78 664 -78 664 5 vdd
rlabel metal1 -76 -116 -76 -116 5 gnd
<< end >>
