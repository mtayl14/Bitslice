magic
tech sky130A
magscale 1 2
timestamp 1701816570
<< nwell >>
rect -98 348 336 706
<< nmos >>
rect 0 -42 30 126
rect 86 -42 116 126
rect 217 0 247 84
<< pmos >>
rect 0 384 30 552
rect 86 384 116 552
rect 217 384 247 552
<< ndiff >>
rect -53 68 0 126
rect -53 16 -45 68
rect -11 16 0 68
rect -53 -42 0 16
rect 30 -42 86 126
rect 116 84 166 126
rect 116 68 217 84
rect 116 16 127 68
rect 206 16 217 68
rect 116 0 217 16
rect 247 68 300 84
rect 247 16 258 68
rect 292 16 300 68
rect 247 0 300 16
rect 116 -42 166 0
<< pdiff >>
rect -53 536 0 552
rect -53 400 -45 536
rect -11 400 0 536
rect -53 384 0 400
rect 30 536 86 552
rect 30 400 41 536
rect 75 400 86 536
rect 30 384 86 400
rect 116 536 217 552
rect 116 400 127 536
rect 206 400 217 536
rect 116 384 217 400
rect 247 536 300 552
rect 247 400 258 536
rect 292 400 300 536
rect 247 384 300 400
<< ndiffc >>
rect -45 16 -11 68
rect 127 16 206 68
rect 258 16 292 68
<< pdiffc >>
rect -45 400 -11 536
rect 41 400 75 536
rect 127 400 206 536
rect 258 400 292 536
<< psubdiff >>
rect -2 -145 23 -111
rect 57 -145 82 -111
rect 136 -145 161 -111
rect 195 -145 220 -111
<< nsubdiff >>
rect 0 636 25 670
rect 59 636 84 670
rect 138 636 163 670
rect 197 636 222 670
<< psubdiffcont >>
rect 23 -145 57 -111
rect 161 -145 195 -111
<< nsubdiffcont >>
rect 25 636 59 670
rect 163 636 197 670
<< poly >>
rect 0 552 30 582
rect 86 552 116 582
rect 217 552 247 582
rect 0 232 30 384
rect -66 216 30 232
rect -66 182 -50 216
rect -16 182 30 216
rect -66 166 30 182
rect 0 126 30 166
rect 86 350 116 384
rect 86 334 175 350
rect 86 300 125 334
rect 159 300 175 334
rect 86 284 175 300
rect 86 126 116 284
rect 217 224 247 384
rect 158 208 247 224
rect 158 174 174 208
rect 208 174 247 208
rect 158 158 247 174
rect 217 84 247 158
rect 217 -30 247 0
rect 0 -72 30 -42
rect 86 -72 116 -42
<< polycont >>
rect -50 182 -16 216
rect 125 300 159 334
rect 174 174 208 208
<< locali >>
rect -98 678 336 697
rect -98 636 25 678
rect 59 636 163 678
rect 197 636 336 678
rect -45 536 -11 636
rect -45 384 -11 400
rect 41 536 75 552
rect -66 216 0 232
rect -66 182 -50 216
rect -16 182 0 216
rect -66 166 0 182
rect 41 192 75 400
rect 127 536 206 636
rect 127 384 206 400
rect 258 536 292 552
rect 109 334 175 350
rect 109 300 125 334
rect 159 300 175 334
rect 109 284 175 300
rect 158 208 224 224
rect 158 192 174 208
rect 41 174 174 192
rect 208 174 224 208
rect 41 158 224 174
rect -45 68 -11 84
rect 41 68 75 158
rect -11 16 75 68
rect 127 68 206 84
rect 258 80 292 400
rect -45 0 -11 16
rect 127 -84 206 16
rect 246 68 304 80
rect 246 16 258 68
rect 292 16 304 68
rect 246 4 304 16
rect 258 0 292 4
rect -100 -92 334 -84
rect -100 -145 23 -92
rect 57 -145 161 -92
rect 195 -145 334 -92
<< viali >>
rect 25 670 59 678
rect 25 644 59 670
rect 163 670 197 678
rect 163 644 197 670
rect -50 182 -16 216
rect 125 300 159 334
rect 258 16 292 68
rect 23 -111 57 -92
rect 23 -126 57 -111
rect 161 -111 195 -92
rect 161 -126 195 -111
<< metal1 >>
rect -98 678 336 697
rect -98 644 25 678
rect 59 644 163 678
rect 197 644 336 678
rect -98 636 336 644
rect 113 340 171 346
rect 113 334 183 340
rect 113 288 125 334
rect 119 282 125 288
rect 177 282 183 334
rect 119 276 183 282
rect -74 234 -10 240
rect -74 182 -68 234
rect -16 228 -10 234
rect -16 182 -4 228
rect -74 176 -4 182
rect -62 170 -4 176
rect 246 74 304 80
rect 246 68 316 74
rect 246 16 258 68
rect 310 16 316 68
rect 246 10 316 16
rect 246 4 304 10
rect -100 -92 334 -84
rect -100 -126 23 -92
rect 57 -126 161 -92
rect 195 -126 334 -92
rect -100 -145 334 -126
<< via1 >>
rect 125 300 159 334
rect 159 300 177 334
rect 125 282 177 300
rect -68 216 -16 234
rect -68 182 -50 216
rect -50 182 -16 216
rect 258 16 292 68
rect 292 16 310 68
<< metal2 >>
rect 119 334 183 340
rect 119 282 125 334
rect 177 282 183 334
rect 119 276 183 282
rect -74 234 -10 240
rect -74 182 -68 234
rect -16 182 -10 234
rect -74 176 -10 182
rect 252 68 316 74
rect 252 16 258 68
rect 310 16 316 68
rect 252 10 316 16
<< labels >>
rlabel via1 284 42 284 42 5 Y
port 3 s
rlabel via1 151 308 151 308 5 B
port 2 s
rlabel via1 -42 208 -42 208 5 A
port 1 s
rlabel polycont 191 191 191 191 5 Y_n
rlabel metal1 -70 -116 -70 -116 5 gnd
rlabel metal1 -70 668 -70 668 5 vdd
<< end >>
