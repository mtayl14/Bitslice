* NGSPICE file created from bitslice.ext - technology: sky130A

.subckt inverter A B gnd vdd
X0 B A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X1 B A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
.ends

.subckt mux21 A B Y S gnd vdd
X0 Y S A vdd sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X1 S_n S gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X2 B S Y gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 S_n S vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
X4 B S_n Y vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.118 ps=1.12 w=0.84 l=0.15
X5 Y S_n A gnd sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.15
.ends

.subckt buffer_fo4 A B gnd vdd
X0 a_n240_0# A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
X1 B a_n240_0# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.47 pd=3.92 as=0.504 ps=3.96 w=1.68 l=0.15
X2 a_n240_0# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X3 vdd a_n240_0# B vdd sky130_fd_pr__pfet_01v8 ad=1.01 pd=7.32 as=0.941 ps=7.28 w=3.36 l=0.15
.ends

.subckt addf A B CI gnd S CO vdd
X0 a_952_521# CI a_870_521# vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.52 as=0.164 ps=1.52 w=1.26 l=0.15
X1 S a_784_115# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.334 pd=3.05 as=0.214 ps=1.6 w=1.26 l=0.15
X2 a_526_115# CI gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X3 a_27_521# B vdd vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X4 a_952_115# CI a_870_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0676 pd=0.78 as=0.0676 ps=0.78 w=0.52 l=0.15
X5 S a_784_115# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.57 as=0.0884 ps=0.86 w=0.52 l=0.15
X6 vdd A a_27_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.334 ps=3.05 w=1.26 l=0.15
X7 a_784_115# CON a_526_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X8 a_27_115# B gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X9 gnd A a_27_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.138 ps=1.57 w=0.52 l=0.15
X10 a_784_115# CON a_526_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X11 CON CI a_27_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X12 vdd A a_368_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.132 ps=1.47 w=1.26 l=0.15
X13 a_526_521# A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X14 CO CON vdd vdd sky130_fd_pr__pfet_01v8 ad=0.334 pd=3.05 as=0.334 ps=3.05 w=1.26 l=0.15
X15 CON CI a_27_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X16 a_870_521# B a_784_115# vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.52 as=0.176 ps=1.54 w=1.26 l=0.15
X17 gnd A a_368_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0546 ps=0.73 w=0.52 l=0.15
X18 a_526_115# A gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X19 CO CON gnd gnd sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.57 as=0.138 ps=1.57 w=0.52 l=0.15
X20 a_870_115# B a_784_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0676 pd=0.78 as=0.0728 ps=0.8 w=0.52 l=0.15
X21 a_368_521# B CON vdd sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.47 as=0.176 ps=1.54 w=1.26 l=0.15
X22 vdd B a_526_521# vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
X23 vdd A a_952_521# vdd sky130_fd_pr__pfet_01v8 ad=0.214 pd=1.6 as=0.164 ps=1.52 w=1.26 l=0.15
X24 a_368_115# B CON gnd sky130_fd_pr__nfet_01v8 ad=0.0546 pd=0.73 as=0.0728 ps=0.8 w=0.52 l=0.15
X25 gnd B a_526_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0728 pd=0.8 as=0.0728 ps=0.8 w=0.52 l=0.15
X26 gnd A a_952_115# gnd sky130_fd_pr__nfet_01v8 ad=0.0884 pd=0.86 as=0.0676 ps=0.78 w=0.52 l=0.15
X27 a_526_521# CI vdd vdd sky130_fd_pr__pfet_01v8 ad=0.176 pd=1.54 as=0.176 ps=1.54 w=1.26 l=0.15
.ends

.subckt d_flip_flop CLK D Q gnd vdd
X0 inverter_1_out common_1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X1 gnd inverter_1_out a_494_0# gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
X2 common_2 CLK_n a_974_426# vdd sky130_fd_pr__pfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 gnd Q a_1248_0# gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
X4 a_974_0# inverter_1_out gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X5 a_220_426# D vdd vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X6 a_494_0# CLK common_1 gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X7 a_1248_0# CLK_n common_2 gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X8 CLK_n CLK vdd vdd sky130_fd_pr__pfet_01v8 ad=0.445 pd=3.89 as=0.445 ps=3.89 w=1.68 l=0.15
X9 common_1 CLK a_220_426# vdd sky130_fd_pr__pfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X10 Q common_2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.34 pd=2.8 as=0.134 ps=1.23 w=0.84 l=0.15
X11 a_1248_426# CLK common_2 vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X12 CLK_n CLK gnd gnd sky130_fd_pr__nfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
X13 common_1 CLK_n a_220_0# gnd sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X14 vdd Q a_1248_426# vdd sky130_fd_pr__pfet_01v8 ad=0.134 pd=1.23 as=0.0819 ps=0.81 w=0.42 l=0.15
X15 common_2 CLK a_974_0# gnd sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X16 inverter_1_out common_1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X17 Q common_2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X18 a_494_426# CLK_n common_1 vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X19 a_974_426# inverter_1_out vdd vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X20 a_220_0# D gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X21 vdd inverter_1_out a_494_426# vdd sky130_fd_pr__pfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
.ends

.subckt and2 A B Y gnd vdd
X0 vdd B Y_n vdd sky130_fd_pr__pfet_01v8 ad=0.212 pd=1.35 as=0.118 ps=1.12 w=0.84 l=0.15
X1 Y Y_n vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.212 ps=1.35 w=0.84 l=0.15
X2 Y Y_n gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.159 ps=1.35 w=0.42 l=0.15
X3 Y_n A vdd vdd sky130_fd_pr__pfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X4 gnd B a_30_n42# gnd sky130_fd_pr__nfet_01v8 ad=0.159 pd=1.35 as=0.118 ps=1.12 w=0.84 l=0.15
X5 a_30_n42# A Y_n gnd sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
.ends

.subckt register D CLK EN Q vdd gnd
Xd_flip_flop_0 and2_0/Y D Q gnd vdd d_flip_flop
Xand2_0 CLK EN and2_0/Y gnd vdd and2
.ends

.subckt bitslice
Xinverter_0 inverter_0/A inverter_0/B VSUBS addf_0/vdd inverter
Xmux21_0 mux21_0/A mux21_0/B mux21_0/Y mux21_0/S VSUBS addf_0/vdd mux21
Xbuffer_fo4_0 buffer_fo4_0/A buffer_fo4_0/B VSUBS addf_0/vdd buffer_fo4
Xaddf_0 addf_0/A addf_0/B addf_0/CI VSUBS addf_0/S addf_0/CO addf_0/vdd addf
Xregister_0 register_0/D register_0/CLK register_0/EN register_0/Q addf_0/vdd VSUBS
+ register
.ends

