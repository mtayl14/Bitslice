magic
tech sky130A
magscale 1 2
timestamp 1701732512
<< nwell >>
rect -98 348 1612 706
<< nmos >>
rect 0 0 30 84
rect 190 0 220 84
rect 298 0 328 84
rect 464 0 494 84
rect 572 0 602 84
rect 680 0 710 84
rect 944 0 974 84
rect 1052 0 1082 84
rect 1218 0 1248 84
rect 1326 0 1356 84
rect 1434 0 1464 84
<< pmos >>
rect 0 384 30 552
rect 190 384 220 552
rect 298 384 328 552
rect 464 384 494 552
rect 572 384 602 552
rect 680 384 710 552
rect 944 384 974 552
rect 1052 384 1082 552
rect 1218 384 1248 552
rect 1326 384 1356 552
rect 1434 384 1464 552
<< ndiff >>
rect -53 68 0 84
rect -53 16 -45 68
rect -11 16 0 68
rect -53 0 0 16
rect 30 68 83 84
rect 30 16 41 68
rect 75 16 83 68
rect 30 0 83 16
rect 137 68 190 84
rect 137 16 145 68
rect 179 16 190 68
rect 137 0 190 16
rect 220 0 298 84
rect 328 68 464 84
rect 328 16 379 68
rect 413 16 464 68
rect 328 0 464 16
rect 494 0 572 84
rect 602 68 680 84
rect 602 16 624 68
rect 658 16 680 68
rect 602 0 680 16
rect 710 68 822 84
rect 710 16 780 68
rect 814 16 822 68
rect 710 0 822 16
rect 891 68 944 84
rect 891 16 899 68
rect 933 16 944 68
rect 891 0 944 16
rect 974 0 1052 84
rect 1082 68 1218 84
rect 1082 16 1133 68
rect 1167 16 1218 68
rect 1082 0 1218 16
rect 1248 0 1326 84
rect 1356 68 1434 84
rect 1356 16 1378 68
rect 1412 16 1434 68
rect 1356 0 1434 16
rect 1464 68 1576 84
rect 1464 16 1534 68
rect 1568 16 1576 68
rect 1464 0 1576 16
<< pdiff >>
rect -53 536 0 552
rect -53 400 -45 536
rect -11 400 0 536
rect -53 384 0 400
rect 30 536 83 552
rect 30 400 41 536
rect 75 400 83 536
rect 30 384 83 400
rect 137 536 190 552
rect 137 400 145 536
rect 179 400 190 536
rect 137 384 190 400
rect 220 384 298 552
rect 328 536 464 552
rect 328 400 379 536
rect 413 400 464 536
rect 328 384 464 400
rect 494 384 572 552
rect 602 536 680 552
rect 602 400 624 536
rect 658 400 680 536
rect 602 384 680 400
rect 710 536 822 552
rect 710 400 780 536
rect 814 400 822 536
rect 710 384 822 400
rect 891 536 944 552
rect 891 400 899 536
rect 933 400 944 536
rect 891 384 944 400
rect 974 384 1052 552
rect 1082 536 1218 552
rect 1082 400 1133 536
rect 1167 400 1218 536
rect 1082 384 1218 400
rect 1248 384 1326 552
rect 1356 536 1434 552
rect 1356 400 1378 536
rect 1412 400 1434 536
rect 1356 384 1434 400
rect 1464 536 1576 552
rect 1464 400 1534 536
rect 1568 400 1576 536
rect 1464 384 1576 400
<< ndiffc >>
rect -45 16 -11 68
rect 41 16 75 68
rect 145 16 179 68
rect 379 16 413 68
rect 624 16 658 68
rect 780 16 814 68
rect 899 16 933 68
rect 1133 16 1167 68
rect 1378 16 1412 68
rect 1534 16 1568 68
<< pdiffc >>
rect -45 400 -11 536
rect 41 400 75 536
rect 145 400 179 536
rect 379 400 413 536
rect 624 400 658 536
rect 780 400 814 536
rect 899 400 933 536
rect 1133 400 1167 536
rect 1378 400 1412 536
rect 1534 400 1568 536
<< psubdiff >>
rect 23 -118 48 -84
rect 82 -118 107 -84
rect 223 -118 248 -84
rect 282 -118 307 -84
rect 423 -118 448 -84
rect 482 -118 507 -84
rect 623 -118 648 -84
rect 682 -118 707 -84
rect 823 -118 848 -84
rect 882 -118 907 -84
rect 1023 -118 1048 -84
rect 1082 -118 1107 -84
rect 1223 -118 1248 -84
rect 1282 -118 1307 -84
rect 1423 -118 1448 -84
rect 1482 -118 1507 -84
<< nsubdiff >>
rect 23 636 48 670
rect 82 636 107 670
rect 223 636 248 670
rect 282 636 307 670
rect 423 636 448 670
rect 482 636 507 670
rect 623 636 648 670
rect 682 636 707 670
rect 823 636 848 670
rect 882 636 907 670
rect 1023 636 1048 670
rect 1082 636 1107 670
rect 1223 636 1248 670
rect 1282 636 1307 670
rect 1423 636 1448 670
rect 1482 636 1507 670
<< psubdiffcont >>
rect 48 -118 82 -84
rect 248 -118 282 -84
rect 448 -118 482 -84
rect 648 -118 682 -84
rect 848 -118 882 -84
rect 1048 -118 1082 -84
rect 1248 -118 1282 -84
rect 1448 -118 1482 -84
<< nsubdiffcont >>
rect 48 636 82 670
rect 248 636 282 670
rect 448 636 482 670
rect 648 636 682 670
rect 848 636 882 670
rect 1048 636 1082 670
rect 1248 636 1282 670
rect 1448 636 1482 670
<< poly >>
rect 0 552 30 582
rect 190 552 220 582
rect 298 552 328 582
rect 464 552 494 582
rect 572 552 602 582
rect 680 552 710 582
rect 944 552 974 582
rect 1052 552 1082 582
rect 1218 552 1248 582
rect 1326 552 1356 582
rect 1434 552 1464 582
rect 0 350 30 384
rect -66 334 30 350
rect -66 300 -50 334
rect -16 300 30 334
rect -66 284 30 300
rect 0 84 30 284
rect 190 252 220 384
rect 298 350 328 384
rect 262 334 328 350
rect 262 300 278 334
rect 312 300 328 334
rect 262 284 328 300
rect 464 350 494 384
rect 464 334 530 350
rect 464 300 480 334
rect 514 300 530 334
rect 464 284 530 300
rect 154 236 220 252
rect 154 202 170 236
rect 204 202 220 236
rect 154 186 220 202
rect 190 84 220 186
rect 572 184 602 384
rect 680 290 710 384
rect 662 274 728 290
rect 662 240 678 274
rect 712 240 728 274
rect 944 250 974 384
rect 1052 350 1082 384
rect 1016 334 1082 350
rect 1016 300 1032 334
rect 1066 300 1082 334
rect 1016 284 1082 300
rect 1218 350 1248 384
rect 1218 334 1284 350
rect 1218 300 1234 334
rect 1268 300 1284 334
rect 1218 284 1284 300
rect 662 224 728 240
rect 878 234 974 250
rect 262 168 328 184
rect 262 134 278 168
rect 312 134 328 168
rect 262 118 328 134
rect 298 84 328 118
rect 464 168 530 184
rect 464 134 480 168
rect 514 134 530 168
rect 464 118 530 134
rect 572 168 638 184
rect 572 134 588 168
rect 622 134 638 168
rect 572 118 638 134
rect 464 84 494 118
rect 572 84 602 118
rect 680 84 710 224
rect 878 200 894 234
rect 928 200 974 234
rect 878 184 974 200
rect 1326 184 1356 384
rect 1434 350 1464 384
rect 1434 334 1500 350
rect 1434 300 1450 334
rect 1484 300 1500 334
rect 1434 284 1500 300
rect 944 84 974 184
rect 1016 168 1082 184
rect 1016 134 1032 168
rect 1066 134 1082 168
rect 1016 118 1082 134
rect 1052 84 1082 118
rect 1218 168 1284 184
rect 1218 134 1234 168
rect 1268 134 1284 168
rect 1218 118 1284 134
rect 1326 168 1392 184
rect 1326 134 1342 168
rect 1376 134 1392 168
rect 1326 118 1392 134
rect 1218 84 1248 118
rect 1326 84 1356 118
rect 1434 84 1464 284
rect 0 -30 30 0
rect 190 -30 220 0
rect 298 -30 328 0
rect 464 -30 494 0
rect 572 -30 602 0
rect 680 -30 710 0
rect 944 -30 974 0
rect 1052 -30 1082 0
rect 1218 -30 1248 0
rect 1326 -30 1356 0
rect 1434 -30 1464 0
<< polycont >>
rect -50 300 -16 334
rect 278 300 312 334
rect 480 300 514 334
rect 170 202 204 236
rect 678 240 712 274
rect 1032 300 1066 334
rect 1234 300 1268 334
rect 278 134 312 168
rect 480 134 514 168
rect 588 134 622 168
rect 894 200 928 234
rect 1450 300 1484 334
rect 1032 134 1066 168
rect 1234 134 1268 168
rect 1342 134 1376 168
<< locali >>
rect -89 670 1578 697
rect -89 636 48 670
rect 82 636 248 670
rect 282 636 448 670
rect 482 636 648 670
rect 682 636 848 670
rect 882 636 1048 670
rect 1082 636 1248 670
rect 1282 636 1448 670
rect 1482 636 1578 670
rect -45 536 -11 636
rect -45 384 -11 400
rect 41 536 75 552
rect -66 334 0 350
rect -66 300 -50 334
rect -16 300 0 334
rect -66 284 0 300
rect 41 152 75 400
rect 145 536 179 636
rect 145 384 179 400
rect 379 536 413 552
rect 262 334 328 350
rect 262 300 278 334
rect 312 300 328 334
rect 262 284 328 300
rect 379 257 413 400
rect 624 536 658 636
rect 624 384 658 400
rect 780 536 814 552
rect 464 334 530 350
rect 464 300 480 334
rect 514 300 530 334
rect 464 284 530 300
rect 662 274 728 290
rect 154 236 220 252
rect 154 202 170 236
rect 204 202 220 236
rect 154 186 220 202
rect 367 245 425 257
rect 367 211 379 245
rect 413 211 425 245
rect 662 240 678 274
rect 712 240 728 274
rect 662 224 728 240
rect 780 234 814 400
rect 899 536 933 636
rect 899 384 933 400
rect 1133 536 1167 552
rect 1016 334 1082 350
rect 1016 300 1032 334
rect 1066 300 1082 334
rect 1016 284 1082 300
rect 878 234 944 250
rect 367 199 425 211
rect 780 200 894 234
rect 928 200 944 234
rect 262 168 328 184
rect 262 152 278 168
rect 41 134 278 152
rect 312 134 328 168
rect 41 118 328 134
rect -45 68 -11 84
rect -45 -84 -11 16
rect 41 68 75 118
rect 41 0 75 16
rect 145 68 179 84
rect 145 -84 179 16
rect 379 68 413 199
rect 379 0 413 16
rect 464 168 530 184
rect 464 134 480 168
rect 514 134 530 168
rect 464 118 530 134
rect 572 168 638 184
rect 572 134 588 168
rect 622 152 638 168
rect 780 152 814 200
rect 878 184 944 200
rect 622 134 814 152
rect 572 118 814 134
rect 1016 168 1082 184
rect 1016 134 1032 168
rect 1066 134 1082 168
rect 1016 118 1082 134
rect 464 22 498 118
rect 624 68 658 84
rect 464 10 522 22
rect 464 -24 476 10
rect 510 -24 522 10
rect 464 -36 522 -24
rect 624 -84 658 16
rect 780 68 814 118
rect 780 0 814 16
rect 899 68 933 84
rect 899 -84 933 16
rect 1133 68 1167 400
rect 1378 536 1412 636
rect 1378 384 1412 400
rect 1534 536 1568 552
rect 1218 334 1284 350
rect 1218 300 1234 334
rect 1268 300 1284 334
rect 1218 284 1284 300
rect 1434 334 1500 350
rect 1434 300 1450 334
rect 1484 300 1500 334
rect 1434 284 1500 300
rect 1218 168 1284 184
rect 1218 134 1234 168
rect 1268 134 1284 168
rect 1218 118 1284 134
rect 1326 168 1392 184
rect 1326 134 1342 168
rect 1376 152 1392 168
rect 1534 152 1568 400
rect 1376 134 1568 152
rect 1326 118 1568 134
rect 1378 68 1412 84
rect 1167 46 1225 58
rect 1167 16 1179 46
rect 1133 12 1179 16
rect 1213 12 1225 46
rect 1133 0 1225 12
rect 1378 -84 1412 16
rect 1534 68 1568 118
rect 1534 0 1568 16
rect -89 -118 48 -84
rect 82 -118 248 -84
rect 282 -118 448 -84
rect 482 -118 648 -84
rect 682 -118 848 -84
rect 882 -118 1048 -84
rect 1082 -118 1248 -84
rect 1282 -118 1448 -84
rect 1482 -118 1578 -84
rect -89 -145 1578 -118
<< viali >>
rect -50 300 -16 334
rect 278 300 312 334
rect 480 300 514 334
rect 170 202 204 236
rect 379 211 413 245
rect 678 240 712 274
rect 1032 300 1066 334
rect 278 134 312 168
rect 480 134 514 168
rect 1032 134 1066 168
rect 476 -24 510 10
rect 1234 300 1268 334
rect 1450 300 1484 334
rect 1234 134 1268 168
rect 1179 12 1213 46
rect 1534 16 1568 50
<< metal1 >>
rect -50 384 1268 418
rect -50 346 -16 384
rect 278 346 312 384
rect 464 346 1066 350
rect 1234 346 1268 384
rect -94 334 -4 346
rect -94 268 -82 334
rect -16 268 -4 334
rect 266 334 324 346
rect 266 300 278 334
rect 312 300 324 334
rect 464 334 1078 346
rect 464 316 480 334
rect 266 288 324 300
rect 468 300 480 316
rect 514 316 1032 334
rect 514 300 526 316
rect 468 288 526 300
rect 1020 300 1032 316
rect 1066 316 1078 334
rect 1222 334 1280 346
rect 1066 308 1128 316
rect 1066 300 1134 308
rect 1020 288 1134 300
rect 1222 300 1234 334
rect 1268 300 1280 334
rect 1222 288 1280 300
rect 1438 334 1496 346
rect 1438 300 1450 334
rect 1484 300 1496 334
rect 1438 288 1496 300
rect -94 256 -4 268
rect 126 268 216 280
rect -50 22 -16 256
rect 126 202 138 268
rect 204 202 216 268
rect 666 274 724 286
rect 126 190 216 202
rect 367 245 425 257
rect 666 245 678 274
rect 367 211 379 245
rect 413 240 678 245
rect 712 240 724 274
rect 413 228 724 240
rect 413 211 711 228
rect 367 199 425 211
rect 266 168 324 180
rect 266 134 278 168
rect 312 134 324 168
rect 266 122 324 134
rect 468 168 526 180
rect 468 134 480 168
rect 514 152 526 168
rect 1020 168 1078 180
rect 1020 152 1032 168
rect 514 134 1032 152
rect 1066 134 1078 168
rect 468 122 1078 134
rect 1106 140 1134 288
rect 1222 168 1280 180
rect 1222 140 1234 168
rect 1106 134 1234 140
rect 1268 134 1280 168
rect 1106 122 1280 134
rect 278 84 312 122
rect 524 118 1064 122
rect 1106 106 1252 122
rect 1106 84 1134 106
rect 278 50 1134 84
rect 1167 56 1225 58
rect 1438 56 1466 288
rect 1528 72 1596 78
rect 1528 62 1534 72
rect 1167 46 1466 56
rect -50 10 522 22
rect -50 -12 476 10
rect 464 -24 476 -12
rect 510 -24 522 10
rect 1167 12 1179 46
rect 1213 22 1466 46
rect 1213 12 1225 22
rect 1167 0 1225 12
rect 1522 16 1534 62
rect 1590 16 1596 72
rect 1522 10 1596 16
rect 1522 4 1580 10
rect 464 -36 522 -24
<< via1 >>
rect -82 300 -50 334
rect -50 300 -16 334
rect -82 268 -16 300
rect 138 236 204 268
rect 138 202 170 236
rect 170 202 204 236
rect 1534 50 1590 72
rect 1534 16 1568 50
rect 1568 16 1590 50
<< metal2 >>
rect -94 334 -4 346
rect -94 268 -82 334
rect -16 268 -4 334
rect -94 256 -4 268
rect 126 268 216 280
rect 126 202 138 268
rect 204 202 216 268
rect 126 190 216 202
rect 1528 72 1596 78
rect 1528 16 1534 72
rect 1590 16 1596 72
rect 1528 10 1596 16
<< labels >>
rlabel metal2 -50 300 -16 334 5 CLK
port 1 s
rlabel metal2 170 202 204 236 5 D
port 2 s
rlabel metal2 1534 16 1590 72 5 Q
port 3 s
rlabel locali -68 -119 -68 -119 5 gnd
rlabel locali -50 670 -50 670 5 vdd
rlabel locali 58 136 58 136 5 CLK_n
rlabel viali 396 228 396 228 5 common_1
rlabel locali 800 218 800 218 5 inverter_1_out
rlabel viali 1196 30 1196 30 5 common_2
<< end >>
