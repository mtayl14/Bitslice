* NGSPICE file created from d_flip_flop.ext - technology: sky130A

.subckt d_flip_flop CLK D Q
X0 gnd inverter_1_out a_494_0# gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
X1 a_220_384# D vdd vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.23 as=0.223 ps=2.21 w=0.84 l=0.15
X2 gnd Q a_1248_0# gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.0819 ps=0.81 w=0.42 l=0.15
X3 CLK_n CLK gnd gnd sky130_fd_pr__nfet_01v8 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.15
X4 common_1 CLK a_220_384# vdd sky130_fd_pr__pfet_01v8 ad=0.286 pd=1.52 as=0.164 ps=1.23 w=0.84 l=0.15
X5 a_974_0# inverter_1_out gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
X6 a_494_0# CLK common_1 gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X7 CLK_n CLK vdd vdd sky130_fd_pr__pfet_01v8 ad=0.223 pd=2.21 as=0.223 ps=2.21 w=0.84 l=0.15
X8 a_1248_0# CLK_n common_2 gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.143 ps=1.1 w=0.42 l=0.15
X9 a_1248_384# CLK common_2 vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.23 as=0.286 ps=1.52 w=0.84 l=0.15
X10 vdd Q a_1248_384# vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.23 as=0.164 ps=1.23 w=0.84 l=0.15
X11 Q common_2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.47 pd=2.8 as=0.164 ps=1.23 w=0.84 l=0.15
X12 common_1 CLK_n a_220_0# gnd sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X13 a_494_384# CLK_n common_1 vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.23 as=0.286 ps=1.52 w=0.84 l=0.15
X14 a_974_384# inverter_1_out vdd vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.23 as=0.223 ps=2.21 w=0.84 l=0.15
X15 common_2 CLK a_974_0# gnd sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.1 as=0.0819 ps=0.81 w=0.42 l=0.15
X16 vdd inverter_1_out a_494_384# vdd sky130_fd_pr__pfet_01v8 ad=0.164 pd=1.23 as=0.164 ps=1.23 w=0.84 l=0.15
X17 inverter_1_out common_1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X18 inverter_1_out common_1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.47 pd=2.8 as=0.164 ps=1.23 w=0.84 l=0.15
X19 common_2 CLK_n a_974_384# vdd sky130_fd_pr__pfet_01v8 ad=0.286 pd=1.52 as=0.164 ps=1.23 w=0.84 l=0.15
X20 Q common_2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.235 pd=1.96 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 a_220_0# D gnd gnd sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.111 ps=1.37 w=0.42 l=0.15
.ends

